* NGSPICE file created from Final2.ext - technology: sky130A

.subckt Dlatch VDD D CLK GND Q NOT_Q
X0 a_430_506# CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=3.24e+12p ps=2.448e+07u w=1e+06u l=150000u
X1 a_94_6# D GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=9e+11p ps=8.6e+06u w=500000u l=150000u
X2 a_1330_6# Q GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=0p ps=0u w=500000u l=150000u
X3 VDD a_480_n20# a_430_506# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Q NOT_Q a_994_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.25e+11p ps=1.5e+06u w=500000u l=150000u
X5 a_994_6# a_94_506# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 a_480_n20# D GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
X7 NOT_Q Q VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_480_n20# D VDD VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X9 VDD CLK a_94_506# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X10 a_430_506# a_480_n20# a_430_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.25e+11p ps=1.5e+06u w=500000u l=150000u
X11 VDD a_430_506# NOT_Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Q a_94_506# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X13 a_94_506# D VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_430_6# CLK GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X15 NOT_Q a_430_506# a_1330_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
X16 VDD NOT_Q Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_94_506# CLK a_94_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
.ends

.subckt inv VDD GND Y A
X0 Y A GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
.ends

.subckt DFF D Q NOT_Q CLK inv_0/GND inv_0/VDD
XDlatch_0 inv_0/VDD D CLK inv_0/GND Dlatch_1/D Dlatch_0/NOT_Q Dlatch
XDlatch_1 inv_0/VDD Dlatch_1/D inv_0/Y inv_0/GND Q NOT_Q Dlatch
Xinv_0 inv_0/VDD inv_0/GND inv_0/Y CLK inv
.ends

.subckt nand2 VDD GND Y A B
X0 a_94_6# A GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=7.2e+11p pd=5.44e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X2 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B a_94_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
.ends

.subckt multiplexor A2 Y2 B2 A3 Y3 B3 A0 Y0 B0 A1 Y1 A6 Y6 B6 A7 Y7 B7 A4 Y4 B4 A5
+ Y5 B5 SEL VDD B1 GND
Xnand2_18 VDD GND nand2_19/A A6 SEL nand2
Xnand2_6 VDD GND nand2_7/A A2 SEL nand2
Xnand2_19 VDD GND Y6 nand2_19/A nand2_21/Y nand2
Xnand2_7 VDD GND Y2 nand2_7/A nand2_8/Y nand2
Xnand2_8 VDD GND nand2_8/Y inv_0/Y B2 nand2
Xnand2_9 VDD GND nand2_9/Y A3 SEL nand2
Xinv_0 VDD GND inv_0/Y SEL inv
Xnand2_20 VDD GND nand2_22/A A7 SEL nand2
Xnand2_21 VDD GND nand2_21/Y inv_0/Y B6 nand2
Xnand2_10 VDD GND Y3 nand2_9/Y nand2_11/Y nand2
Xnand2_22 VDD GND Y7 nand2_22/A nand2_23/Y nand2
Xnand2_11 VDD GND nand2_11/Y inv_0/Y B3 nand2
Xnand2_23 VDD GND nand2_23/Y inv_0/Y B7 nand2
Xnand2_12 VDD GND nand2_13/A A4 SEL nand2
Xnand2_0 VDD GND nand2_1/A A0 SEL nand2
Xnand2_13 VDD GND Y4 nand2_13/A nand2_14/Y nand2
Xnand2_2 VDD GND nand2_2/Y inv_0/Y B0 nand2
Xnand2_1 VDD GND Y0 nand2_1/A nand2_2/Y nand2
Xnand2_14 VDD GND nand2_14/Y inv_0/Y B4 nand2
Xnand2_3 VDD GND nand2_4/B inv_0/Y B1 nand2
Xnand2_16 VDD GND Y5 nand2_16/A nand2_17/Y nand2
Xnand2_15 VDD GND nand2_16/A A5 SEL nand2
Xnand2_4 VDD GND Y1 nand2_5/Y nand2_4/B nand2
Xnand2_17 VDD GND nand2_17/Y inv_0/Y B5 nand2
Xnand2_5 VDD GND nand2_5/Y A1 SEL nand2
.ends

*.subckt Final2 CLK A B Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
XDFF_0 DFF_0/D DFF_0/Q DFF_0/D CLK GND VDD DFF
XDFF_1 DFF_1/D DFF_1/Q DFF_1/D DFF_0/Q GND VDD DFF
XDFF_3 DFF_3/D DFF_3/Q DFF_3/D DFF_1/Q GND VDD DFF
XDFF_2 DFF_2/D DFF_2/Q DFF_2/D DFF_3/Q GND VDD DFF
Xmultiplexor_0 multiplexor_1/Y2 multiplexor_2/B2 DFF_2/Q multiplexor_1/Y3 multiplexor_2/B3
+ multiplexor_1/A4 multiplexor_1/Y0 multiplexor_2/B0 DFF_1/Q multiplexor_1/Y1 multiplexor_2/B1
+ multiplexor_1/Y6 multiplexor_2/B6 DFF_7/Q multiplexor_1/Y7 multiplexor_2/B7 DFF_8/Q
+ multiplexor_1/Y4 multiplexor_2/B4 DFF_4/Q multiplexor_1/Y5 multiplexor_2/B5 DFF_6/Q
+ B VDD DFF_3/Q GND multiplexor
XDFF_4 DFF_4/D DFF_4/Q DFF_4/D DFF_5/Q GND VDD DFF
Xmultiplexor_1 DFF_3/Q multiplexor_1/Y2 DFF_3/D DFF_2/Q multiplexor_1/Y3 DFF_2/D DFF_0/Q
+ multiplexor_1/Y0 DFF_0/D DFF_1/Q multiplexor_1/Y1 DFF_6/Q multiplexor_1/Y6 DFF_6/D
+ DFF_7/Q multiplexor_1/Y7 DFF_7/D multiplexor_1/A4 multiplexor_1/Y4 DFF_5/D DFF_4/Q
+ multiplexor_1/Y5 DFF_4/D DFF_8/D VDD DFF_1/D GND multiplexor
XDFF_5 DFF_5/D DFF_5/Q DFF_5/D DFF_2/Q GND VDD DFF
Xmultiplexor_2 DFF_8/Q Y2 multiplexor_2/B2 DFF_8/Q Y3 multiplexor_2/B3 DFF_8/Q Y0
+ multiplexor_2/B0 DFF_8/Q Y1 DFF_8/Q Y6 multiplexor_2/B6 DFF_8/Q Y7 multiplexor_2/B7
+ DFF_8/Q Y4 multiplexor_2/B4 DFF_8/Q Y5 multiplexor_2/B5 A VDD multiplexor_2/B1 GND
+ multiplexor
XDFF_6 DFF_6/D DFF_6/Q DFF_6/D DFF_4/Q GND VDD DFF
XDFF_7 DFF_7/D DFF_7/Q DFF_7/D DFF_6/Q GND VDD DFF
XDFF_8 DFF_8/D DFF_8/Q DFF_8/D DFF_7/Q GND VDD DFF
*.ends

