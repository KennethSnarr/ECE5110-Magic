* NGSPICE file created from 9bit_count.ext - technology: sky130A

.subckt Dlatch VDD D CLK GND Q NOT_Q
X0 a_430_506# CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=3.24e+12p ps=2.448e+07u w=1e+06u l=150000u
X1 a_94_6# D GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=9e+11p ps=8.6e+06u w=500000u l=150000u
X2 a_1330_6# Q GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=0p ps=0u w=500000u l=150000u
X3 VDD a_480_n20# a_430_506# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Q NOT_Q a_994_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.25e+11p ps=1.5e+06u w=500000u l=150000u
X5 a_994_6# a_94_506# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 a_480_n20# D GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
X7 NOT_Q Q VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_480_n20# D VDD VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X9 VDD CLK a_94_506# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X10 a_430_506# a_480_n20# a_430_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.25e+11p ps=1.5e+06u w=500000u l=150000u
X11 VDD a_430_506# NOT_Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Q a_94_506# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X13 a_94_506# D VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_430_6# CLK GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X15 NOT_Q a_430_506# a_1330_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
X16 VDD NOT_Q Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_94_506# CLK a_94_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
.ends

.subckt inv VDD GND Y A
X0 Y A GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
.ends

.subckt DFF D Q NOT_Q CLK inv_0/GND inv_0/VDD
XDlatch_0 inv_0/VDD D CLK inv_0/GND Dlatch_1/D Dlatch_0/NOT_Q Dlatch
XDlatch_1 inv_0/VDD Dlatch_1/D inv_0/Y inv_0/GND Q NOT_Q Dlatch
Xinv_0 inv_0/VDD inv_0/GND inv_0/Y CLK inv
.ends

*.subckt x9bit_count CLK Y
XDFF_0 DFF_0/D DFF_0/Q DFF_0/D DFF_8/Q GND VDD DFF
XDFF_1 DFF_1/D DFF_1/Q DFF_1/D DFF_0/Q GND VDD DFF
XDFF_2 DFF_2/D DFF_2/Q DFF_2/D DFF_1/Q GND VDD DFF
XDFF_3 DFF_3/D DFF_3/Q DFF_3/D DFF_2/Q GND VDD DFF
XDFF_4 DFF_4/D Y DFF_4/NOT_Q DFF_5/Q GND VDD DFF
XDFF_5 DFF_5/D DFF_5/Q DFF_5/D DFF_6/Q GND VDD DFF
XDFF_6 DFF_6/D DFF_6/Q DFF_6/D DFF_7/Q GND VDD DFF
XDFF_7 DFF_7/D DFF_7/Q DFF_7/D DFF_3/Q GND VDD DFF
XDFF_8 DFF_8/D DFF_8/Q DFF_8/D CLK GND VDD DFF
*.ends

