* NGSPICE file created from nor2.ext - technology: sky130A

*.subckt nor2 VDD GND Y A B
X0 Y A GND GND sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.78e+06u as=3.6e+11p ps=3.44e+06u w=500000u l=150000u
X1 GND B Y GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2 Y B a_94_506# VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=2.5e+11p ps=2.5e+06u w=1e+06u l=150000u
X3 a_94_506# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
*.ends

