magic
tech sky130A
magscale 1 2
timestamp 1680222599
<< poly >>
rect 1716 104 1746 106
<< locali >>
rect -264 864 3840 960
rect -186 433 -159 464
rect -125 433 -120 464
rect -84 312 -18 630
rect 400 528 466 562
rect 400 494 412 528
rect 446 494 466 528
rect 38 380 70 446
rect 400 432 466 494
rect 640 449 706 464
rect 640 434 657 449
rect 190 414 256 432
rect 190 380 203 414
rect 237 380 256 414
rect 640 398 650 434
rect 691 415 706 449
rect 690 398 706 415
rect 190 366 256 380
rect 394 359 460 390
rect -84 278 -74 312
rect -40 278 -18 312
rect -84 230 -18 278
rect 532 270 598 302
rect 742 323 808 630
rect 908 449 974 464
rect 908 415 921 449
rect 955 415 974 449
rect 908 398 974 415
rect 1010 449 1076 630
rect 1112 480 1178 512
rect 1010 415 1022 449
rect 1056 415 1076 449
rect 1010 328 1076 415
rect 1308 398 1340 464
rect 1376 448 1442 630
rect 1376 414 1387 448
rect 1421 414 1442 448
rect 742 289 759 323
rect 793 289 808 323
rect 742 230 808 289
rect 1376 230 1442 414
rect 1576 398 1608 464
rect 1644 461 1710 542
rect 1644 427 1658 461
rect 1692 427 1710 461
rect 1644 230 1710 427
rect 1904 398 1970 422
rect 1746 316 1774 382
rect 2006 230 2072 630
rect 2144 398 2210 424
rect 2246 366 2312 630
rect 2514 555 2580 630
rect 2514 521 2525 555
rect 2559 521 2580 555
rect 2412 398 2444 464
rect 2246 332 2263 366
rect 2297 332 2312 366
rect 2246 230 2312 332
rect 2514 328 2580 521
rect 2774 398 2802 464
rect 2876 317 2942 630
rect 2998 427 3064 446
rect 3360 432 3426 562
rect 3600 447 3666 464
rect 2998 393 3013 427
rect 3047 393 3064 427
rect 2998 380 3064 393
rect 3600 413 3606 447
rect 3640 413 3666 447
rect 3600 398 3666 413
rect 2876 283 2887 317
rect 2921 283 2942 317
rect 2876 230 2942 283
rect 3702 330 3768 630
rect 3751 276 3768 330
rect 3702 230 3768 276
rect -264 0 3840 96
<< viali >>
rect -159 433 -125 466
rect -186 398 -120 433
rect 412 494 446 528
rect 70 380 104 446
rect 657 434 691 449
rect 203 380 237 414
rect 650 415 691 434
rect 650 394 690 415
rect 394 324 460 359
rect -74 278 -40 312
rect 532 302 598 336
rect 921 415 955 449
rect 1112 512 1178 546
rect 1022 415 1056 449
rect 1274 398 1308 464
rect 1387 414 1421 448
rect 759 289 793 323
rect 1542 398 1576 464
rect 1658 427 1692 461
rect 1904 422 1970 464
rect 1774 316 1812 382
rect 2144 424 2210 464
rect 2525 521 2559 555
rect 2444 398 2478 464
rect 2263 332 2297 366
rect 2616 480 2682 546
rect 2802 398 2840 464
rect 3013 393 3047 427
rect 3150 366 3216 432
rect 3606 413 3640 447
rect 3354 324 3420 390
rect 2887 283 2921 317
rect 3492 270 3558 336
rect 3697 276 3751 330
<< metal1 >>
rect 407 618 3645 661
rect -157 520 235 551
rect 407 540 450 618
rect 2513 558 2571 561
rect 2157 555 2571 558
rect 1100 546 1190 552
rect -157 472 -126 520
rect -171 466 -113 472
rect -171 439 -159 466
rect -198 433 -159 439
rect -125 439 -113 466
rect 64 452 110 458
rect -125 433 -108 439
rect -198 398 -186 433
rect -120 398 -108 433
rect -198 392 -108 398
rect -170 140 -135 392
rect 55 374 61 452
rect 113 374 119 452
rect 204 426 235 520
rect 406 528 452 540
rect 406 494 412 528
rect 446 494 452 528
rect 406 482 452 494
rect 657 512 1112 546
rect 1178 512 1190 546
rect 657 461 691 512
rect 1100 506 1190 512
rect 2157 521 2525 555
rect 2559 521 2571 555
rect 2617 552 2682 618
rect 2157 518 2571 521
rect 1268 464 1314 476
rect 651 449 697 461
rect 651 446 657 449
rect 644 440 657 446
rect 691 440 697 449
rect 197 414 243 426
rect 197 380 203 414
rect 237 380 243 414
rect 64 368 110 374
rect 197 368 243 380
rect 290 407 582 440
rect -86 312 -28 318
rect -86 278 -74 312
rect -40 311 -28 312
rect 290 311 323 407
rect 382 359 472 365
rect 382 324 394 359
rect 460 324 472 359
rect 549 342 582 407
rect 696 403 697 440
rect 915 449 961 461
rect 915 415 921 449
rect 955 415 961 449
rect 915 403 961 415
rect 1010 449 1068 455
rect 1010 415 1022 449
rect 1056 448 1068 449
rect 1268 448 1274 464
rect 1056 415 1274 448
rect 1010 409 1068 415
rect 644 382 696 388
rect 382 318 472 324
rect 520 336 610 342
rect -40 278 323 311
rect -86 272 -28 278
rect 410 220 445 318
rect 520 302 532 336
rect 598 302 610 336
rect 520 296 610 302
rect 753 323 799 335
rect 753 289 759 323
rect 793 289 799 323
rect 753 277 799 289
rect 758 220 793 277
rect 410 185 793 220
rect 920 140 955 403
rect 1268 398 1274 415
rect 1308 398 1314 464
rect 1536 464 1582 476
rect 2157 470 2197 518
rect 2513 515 2571 518
rect 2604 546 2694 552
rect 2604 480 2616 546
rect 2682 480 2694 546
rect 1375 448 1433 454
rect 1375 414 1387 448
rect 1421 447 1433 448
rect 1536 447 1542 464
rect 1421 415 1542 447
rect 1421 414 1433 415
rect 1375 408 1433 414
rect 1268 386 1314 398
rect 1536 398 1542 415
rect 1576 398 1582 464
rect 1646 465 1704 467
rect 1892 465 1982 470
rect 1646 464 1982 465
rect 1646 461 1904 464
rect 1646 427 1658 461
rect 1692 427 1904 461
rect 1646 422 1904 427
rect 1970 422 1982 464
rect 1646 421 1704 422
rect 1892 416 1982 422
rect 2132 464 2222 470
rect 2132 424 2144 464
rect 2210 424 2222 464
rect 2132 418 2222 424
rect 2438 464 2484 476
rect 2604 474 2694 480
rect 1536 386 1582 398
rect 2438 398 2444 464
rect 2478 411 2484 464
rect 2796 464 2846 476
rect 2796 411 2802 464
rect 2478 398 2802 411
rect 2840 450 2846 464
rect 2840 439 3049 450
rect 3162 444 3205 618
rect 3607 459 3639 618
rect 3600 447 3646 459
rect 2840 427 3053 439
rect 2840 412 3013 427
rect 2840 398 2846 412
rect 1768 382 1818 394
rect 2438 386 2846 398
rect 3007 393 3013 412
rect 3047 393 3053 427
rect 1768 316 1774 382
rect 1812 368 1818 382
rect 2444 377 2841 386
rect 3007 381 3053 393
rect 3144 432 3222 444
rect 2251 368 2309 372
rect 1812 366 2309 368
rect 1812 332 2263 366
rect 2297 332 2309 366
rect 3144 366 3150 432
rect 3216 366 3222 432
rect 3600 413 3606 447
rect 3640 413 3646 447
rect 3600 401 3646 413
rect 3144 354 3222 366
rect 3342 390 3432 396
rect 1812 330 2309 332
rect 1812 316 1818 330
rect 2251 326 2309 330
rect 3342 324 3354 390
rect 3420 324 3432 390
rect 1768 304 1818 316
rect 2875 322 2933 323
rect 3342 322 3432 324
rect 2875 318 3432 322
rect 3486 336 3564 348
rect 2875 317 3409 318
rect 2875 283 2887 317
rect 2921 283 3409 317
rect 2875 278 3409 283
rect 2875 277 2933 278
rect 3486 270 3492 336
rect 3558 330 3763 336
rect 3558 276 3697 330
rect 3751 276 3763 330
rect 3558 270 3763 276
rect 3486 258 3564 270
rect -170 105 955 140
<< via1 >>
rect 61 446 113 452
rect 61 380 70 446
rect 70 380 104 446
rect 104 380 113 446
rect 61 374 113 380
rect 644 434 657 440
rect 657 434 691 440
rect 644 394 650 434
rect 650 415 691 434
rect 691 415 696 440
rect 650 394 690 415
rect 690 394 696 415
rect 644 388 696 394
<< metal2 >>
rect 61 452 113 458
rect 638 428 644 440
rect 113 399 644 428
rect 638 388 644 399
rect 696 388 702 440
rect 61 368 113 374
use inv  inv_0
timestamp 1679616770
transform 1 0 642 0 1 124
box -84 -124 242 852
use inv  inv_1
timestamp 1679616770
transform 1 0 -184 0 1 124
box -84 -124 242 852
use inv  inv_2
timestamp 1679616770
transform 1 0 1276 0 1 124
box -84 -124 242 852
use inv  inv_3
timestamp 1679616770
transform 1 0 1906 0 1 124
box -84 -124 242 852
use inv  inv_4
timestamp 1679616770
transform 1 0 2146 0 1 124
box -84 -124 242 852
use inv  inv_5
timestamp 1679616770
transform 1 0 2776 0 1 124
box -84 -124 242 852
use inv  inv_6
timestamp 1679616770
transform 1 0 3602 0 1 124
box -84 -124 242 852
use nand2  nand2_0
timestamp 1676660346
transform 1 0 910 0 1 124
box -84 -124 350 852
use nand2  nand2_1
timestamp 1676660346
transform 1 0 2414 0 1 124
box -84 -124 350 852
use nor2  nor2_0
timestamp 1676660012
transform 1 0 1544 0 1 124
box -84 -124 350 852
use xor2  xor2_0
timestamp 1677800174
transform 1 0 84 0 1 124
box -84 -124 566 852
use xor2  xor2_1
timestamp 1677800174
transform 1 0 3044 0 1 124
box -84 -124 566 852
<< labels >>
flabel locali s 3360 432 3426 562 0 FreeSerif 320 0 0 0 S
port 0 nsew
flabel locali s 2998 380 3064 446 0 FreeSerif 320 0 0 0 C_in
port 7 nsew
flabel locali s 2006 230 2072 630 0 FreeSerif 320 0 0 0 C_out
port 10 nsew
flabel locali s -186 398 -120 464 0 FreeSerif 320 0 0 0 A
port 1 nsew
flabel locali s 640 398 706 464 0 FreeSerif 320 0 0 0 B
port 2 nsew
<< end >>
