* NGSPICE file created from DFF.ext - technology: sky130A

*.subckt DFF VDD D CLK GND Q NOT_Q
X0 a_430_506# CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=3.24e+12p ps=2.448e+07u w=1e+06u l=150000u
X1 a_94_6# D GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=9e+11p ps=8.6e+06u w=500000u l=150000u
X2 a_1330_6# Q GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=0p ps=0u w=500000u l=150000u
X3 VDD a_480_n20# a_430_506# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Q NOT_Q a_994_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.25e+11p ps=1.5e+06u w=500000u l=150000u
X5 a_994_6# a_94_506# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 a_480_n20# D GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
X7 NOT_Q Q VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_480_n20# D VDD VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=0p ps=0u w=1e+06u l=150000u
X9 VDD CLK a_94_506# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X10 a_430_506# a_480_n20# a_430_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.25e+11p ps=1.5e+06u w=500000u l=150000u
X11 VDD a_430_506# NOT_Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Q a_94_506# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X13 a_94_506# D VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_430_6# CLK GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X15 NOT_Q a_430_506# a_1330_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
X16 VDD NOT_Q Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_94_506# CLK a_94_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
*.ends

