magic
tech sky130A
timestamp 1676660346
<< nwell >>
rect -42 135 175 426
<< nmos >>
rect 32 3 47 53
rect 72 3 87 53
<< pmos >>
rect 32 253 47 353
rect 86 253 101 353
<< ndiff >>
rect -4 45 32 53
rect -4 11 4 45
rect 21 11 32 45
rect -4 3 32 11
rect 47 3 72 53
rect 87 45 123 53
rect 87 11 98 45
rect 115 11 123 45
rect 87 3 123 11
<< pdiff >>
rect -4 345 32 353
rect -4 261 4 345
rect 21 261 32 345
rect -4 253 32 261
rect 47 345 86 353
rect 47 261 58 345
rect 75 261 86 345
rect 47 253 86 261
rect 101 345 137 353
rect 101 261 112 345
rect 129 261 137 345
rect 101 253 137 261
<< ndiffc >>
rect 4 11 21 45
rect 98 11 115 45
<< pdiffc >>
rect 4 261 21 345
rect 58 261 75 345
rect 112 261 129 345
<< psubdiff >>
rect -4 -52 8 -24
rect 111 -52 123 -24
<< nsubdiff >>
rect 3 380 15 408
rect 118 380 130 408
<< psubdiffcont >>
rect 8 -52 111 -24
<< nsubdiffcont >>
rect 15 380 118 408
<< poly >>
rect 32 353 47 366
rect 86 353 101 366
rect 32 170 47 253
rect -1 162 47 170
rect -1 145 7 162
rect 24 145 47 162
rect -1 137 47 145
rect 32 53 47 137
rect 86 211 101 253
rect 86 203 134 211
rect 86 186 109 203
rect 126 186 134 203
rect 86 178 134 186
rect 86 99 101 178
rect 72 84 101 99
rect 72 53 87 84
rect 32 -10 47 3
rect 72 -10 87 3
<< polycont >>
rect 7 145 24 162
rect 109 186 126 203
<< locali >>
rect -40 408 173 418
rect -40 380 15 408
rect 118 380 173 408
rect -40 370 173 380
rect -4 345 29 370
rect -4 261 4 345
rect 21 261 29 345
rect -4 253 29 261
rect 50 345 83 353
rect 50 261 58 345
rect 75 261 83 345
rect -1 162 32 170
rect -1 145 7 162
rect 24 145 32 162
rect -1 137 32 145
rect 50 135 83 261
rect 104 345 137 370
rect 104 261 112 345
rect 129 261 137 345
rect 104 253 137 261
rect 101 203 134 211
rect 101 186 109 203
rect 126 186 134 203
rect 101 178 134 186
rect 50 102 123 135
rect -4 45 29 53
rect -4 11 4 45
rect 21 11 29 45
rect -4 -14 29 11
rect 90 45 123 102
rect 90 11 98 45
rect 115 11 123 45
rect 90 3 123 11
rect -40 -24 173 -14
rect -40 -52 8 -24
rect 111 -52 173 -24
rect -40 -62 173 -52
<< labels >>
flabel locali -1 137 32 170 0 FreeSerif 80 0 0 0 A
port 3 nsew
flabel locali 101 178 134 211 0 FreeSerif 80 0 0 0 B
port 8 nsew
flabel locali 50 102 83 253 0 FreeSerif 80 0 0 0 Y
port 2 nsew
flabel locali -40 370 173 418 0 FreeSerif 80 0 0 0 VDD!
port 0 nsew
flabel locali -40 -62 173 -14 0 FreeSerif 80 0 0 0 GND!
port 1 nsew
<< end >>
