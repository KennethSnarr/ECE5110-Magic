* NGSPICE file created from full_adder.ext - technology: sky130A

.subckt nor2 VDD GND Y A B
X0 Y A GND GND sky130_fd_pr__nfet_01v8 ad=1.95e+11p pd=1.78e+06u as=3.6e+11p ps=3.44e+06u w=500000u l=150000u
X1 GND B Y GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X2 Y B a_94_506# VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=2.5e+11p ps=2.5e+06u w=1e+06u l=150000u
X3 a_94_506# A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
.ends

.subckt xor2 VDD GND Y A B NOT_A NOT_B
X0 a_94_6# B GND GND sky130_fd_pr__nfet_01v8 ad=1.05e+11p pd=1.42e+06u as=3.9e+11p ps=3.56e+06u w=500000u l=150000u
X1 a_274_6# NOT_B Y GND sky130_fd_pr__nfet_01v8 ad=1.05e+11p pd=1.42e+06u as=1.95e+11p ps=1.78e+06u w=500000u l=150000u
X2 Y A a_94_6# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X3 a_n8_438# A VDD VDD sky130_fd_pr__pfet_01v8 ad=1.14e+12p pd=8.28e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X4 Y NOT_B a_n8_438# VDD sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u l=150000u
X5 GND NOT_A a_274_6# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=150000u
X6 a_n8_438# NOT_A Y VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VDD B a_n8_438# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt inv VDD GND Y A
X0 Y A GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
.ends

.subckt nand2 VDD GND Y A B
X0 a_94_6# A GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=7.2e+11p pd=5.44e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X2 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B a_94_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
.ends

.subckt half_adder S A B C_out GND VDD
Xxor2_0 VDD GND S A B inv_2/Y inv_1/Y xor2
Xinv_0 VDD GND C_out inv_0/A inv
Xinv_1 VDD GND inv_1/Y B inv
Xinv_2 VDD GND inv_2/Y A inv
Xnand2_0 VDD GND inv_0/A A B nand2
.ends

*.subckt full_adder S A B C_out
Xnor2_0 inv_0/VDD inv_0/GND inv_0/A nor2_0/A nor2_0/B nor2
Xhalf_adder_0 half_adder_1/A A B nor2_0/A inv_0/GND inv_0/VDD half_adder
Xhalf_adder_1 S half_adder_1/A half_adder_1/B nor2_0/B inv_0/GND inv_0/VDD half_adder
Xinv_0 inv_0/VDD inv_0/GND C_out inv_0/A inv
*.ends

