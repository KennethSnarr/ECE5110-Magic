magic
tech sky130A
magscale 1 2
timestamp 1681156228
<< nwell >>
rect 0 848 13866 1430
<< nmos >>
rect 148 1594 178 1694
rect 416 1594 446 1694
rect 496 1594 526 1694
rect 752 1594 782 1694
rect 832 1594 862 1694
rect 1088 1594 1118 1694
rect 1316 1594 1346 1694
rect 1396 1594 1426 1694
rect 1652 1594 1682 1694
rect 1732 1594 1762 1694
rect 1988 1594 2018 1694
rect 2068 1594 2098 1694
rect 2324 1594 2354 1694
rect 2404 1594 2434 1694
rect 2660 1594 2690 1694
rect 2888 1594 2918 1694
rect 2968 1594 2998 1694
rect 3224 1594 3254 1694
rect 3304 1594 3334 1694
rect 3600 1594 3630 1694
rect 3868 1594 3898 1694
rect 3948 1594 3978 1694
rect 4204 1594 4234 1694
rect 4284 1594 4314 1694
rect 4540 1594 4570 1694
rect 4768 1594 4798 1694
rect 4848 1594 4878 1694
rect 5104 1594 5134 1694
rect 5184 1594 5214 1694
rect 5440 1594 5470 1694
rect 5520 1594 5550 1694
rect 5776 1594 5806 1694
rect 5856 1594 5886 1694
rect 6112 1594 6142 1694
rect 6340 1594 6370 1694
rect 6420 1594 6450 1694
rect 6676 1594 6706 1694
rect 6756 1594 6786 1694
rect 7052 1594 7082 1694
rect 7320 1594 7350 1694
rect 7400 1594 7430 1694
rect 7656 1594 7686 1694
rect 7736 1594 7766 1694
rect 7992 1594 8022 1694
rect 8220 1594 8250 1694
rect 8300 1594 8330 1694
rect 8556 1594 8586 1694
rect 8636 1594 8666 1694
rect 8892 1594 8922 1694
rect 8972 1594 9002 1694
rect 9228 1594 9258 1694
rect 9308 1594 9338 1694
rect 9564 1594 9594 1694
rect 9792 1594 9822 1694
rect 9872 1594 9902 1694
rect 10128 1594 10158 1694
rect 10208 1594 10238 1694
rect 10504 1594 10534 1694
rect 10772 1594 10802 1694
rect 10852 1594 10882 1694
rect 11108 1594 11138 1694
rect 11188 1594 11218 1694
rect 11444 1594 11474 1694
rect 11672 1594 11702 1694
rect 11752 1594 11782 1694
rect 12008 1594 12038 1694
rect 12088 1594 12118 1694
rect 12344 1594 12374 1694
rect 12424 1594 12454 1694
rect 12680 1594 12710 1694
rect 12760 1594 12790 1694
rect 13016 1594 13046 1694
rect 13244 1594 13274 1694
rect 13324 1594 13354 1694
rect 13580 1594 13610 1694
rect 13660 1594 13690 1694
<< pmos >>
rect 148 994 178 1194
rect 416 994 446 1194
rect 524 994 554 1194
rect 752 994 782 1194
rect 860 994 890 1194
rect 1088 994 1118 1194
rect 1316 994 1346 1194
rect 1424 994 1454 1194
rect 1652 994 1682 1194
rect 1760 994 1790 1194
rect 1988 994 2018 1194
rect 2096 994 2126 1194
rect 2324 994 2354 1194
rect 2432 994 2462 1194
rect 2660 994 2690 1194
rect 2888 994 2918 1194
rect 2996 994 3026 1194
rect 3224 994 3254 1194
rect 3332 994 3362 1194
rect 3600 994 3630 1194
rect 3868 994 3898 1194
rect 3976 994 4006 1194
rect 4204 994 4234 1194
rect 4312 994 4342 1194
rect 4540 994 4570 1194
rect 4768 994 4798 1194
rect 4876 994 4906 1194
rect 5104 994 5134 1194
rect 5212 994 5242 1194
rect 5440 994 5470 1194
rect 5548 994 5578 1194
rect 5776 994 5806 1194
rect 5884 994 5914 1194
rect 6112 994 6142 1194
rect 6340 994 6370 1194
rect 6448 994 6478 1194
rect 6676 994 6706 1194
rect 6784 994 6814 1194
rect 7052 994 7082 1194
rect 7320 994 7350 1194
rect 7428 994 7458 1194
rect 7656 994 7686 1194
rect 7764 994 7794 1194
rect 7992 994 8022 1194
rect 8220 994 8250 1194
rect 8328 994 8358 1194
rect 8556 994 8586 1194
rect 8664 994 8694 1194
rect 8892 994 8922 1194
rect 9000 994 9030 1194
rect 9228 994 9258 1194
rect 9336 994 9366 1194
rect 9564 994 9594 1194
rect 9792 994 9822 1194
rect 9900 994 9930 1194
rect 10128 994 10158 1194
rect 10236 994 10266 1194
rect 10504 994 10534 1194
rect 10772 994 10802 1194
rect 10880 994 10910 1194
rect 11108 994 11138 1194
rect 11216 994 11246 1194
rect 11444 994 11474 1194
rect 11672 994 11702 1194
rect 11780 994 11810 1194
rect 12008 994 12038 1194
rect 12116 994 12146 1194
rect 12344 994 12374 1194
rect 12452 994 12482 1194
rect 12680 994 12710 1194
rect 12788 994 12818 1194
rect 13016 994 13046 1194
rect 13244 994 13274 1194
rect 13352 994 13382 1194
rect 13580 994 13610 1194
rect 13688 994 13718 1194
<< ndiff >>
rect 76 1678 148 1694
rect 76 1610 92 1678
rect 126 1610 148 1678
rect 76 1594 148 1610
rect 178 1678 250 1694
rect 178 1610 200 1678
rect 234 1610 250 1678
rect 178 1594 250 1610
rect 344 1678 416 1694
rect 344 1610 360 1678
rect 394 1610 416 1678
rect 344 1594 416 1610
rect 446 1594 496 1694
rect 526 1678 598 1694
rect 526 1610 548 1678
rect 582 1610 598 1678
rect 526 1594 598 1610
rect 680 1678 752 1694
rect 680 1610 696 1678
rect 730 1610 752 1678
rect 680 1594 752 1610
rect 782 1594 832 1694
rect 862 1678 934 1694
rect 862 1610 884 1678
rect 918 1610 934 1678
rect 862 1594 934 1610
rect 1016 1678 1088 1694
rect 1016 1610 1032 1678
rect 1066 1610 1088 1678
rect 1016 1594 1088 1610
rect 1118 1678 1190 1694
rect 1118 1610 1140 1678
rect 1174 1610 1190 1678
rect 1118 1594 1190 1610
rect 1244 1678 1316 1694
rect 1244 1610 1260 1678
rect 1294 1610 1316 1678
rect 1244 1594 1316 1610
rect 1346 1594 1396 1694
rect 1426 1678 1498 1694
rect 1426 1610 1448 1678
rect 1482 1610 1498 1678
rect 1426 1594 1498 1610
rect 1580 1678 1652 1694
rect 1580 1610 1596 1678
rect 1630 1610 1652 1678
rect 1580 1594 1652 1610
rect 1682 1594 1732 1694
rect 1762 1678 1834 1694
rect 1762 1610 1784 1678
rect 1818 1610 1834 1678
rect 1762 1594 1834 1610
rect 1916 1678 1988 1694
rect 1916 1610 1932 1678
rect 1966 1610 1988 1678
rect 1916 1594 1988 1610
rect 2018 1594 2068 1694
rect 2098 1678 2170 1694
rect 2098 1610 2120 1678
rect 2154 1610 2170 1678
rect 2098 1594 2170 1610
rect 2252 1678 2324 1694
rect 2252 1610 2268 1678
rect 2302 1610 2324 1678
rect 2252 1594 2324 1610
rect 2354 1594 2404 1694
rect 2434 1678 2506 1694
rect 2434 1610 2456 1678
rect 2490 1610 2506 1678
rect 2434 1594 2506 1610
rect 2588 1678 2660 1694
rect 2588 1610 2604 1678
rect 2638 1610 2660 1678
rect 2588 1594 2660 1610
rect 2690 1678 2762 1694
rect 2690 1610 2712 1678
rect 2746 1610 2762 1678
rect 2690 1594 2762 1610
rect 2816 1678 2888 1694
rect 2816 1610 2832 1678
rect 2866 1610 2888 1678
rect 2816 1594 2888 1610
rect 2918 1594 2968 1694
rect 2998 1678 3070 1694
rect 2998 1610 3020 1678
rect 3054 1610 3070 1678
rect 2998 1594 3070 1610
rect 3152 1678 3224 1694
rect 3152 1610 3168 1678
rect 3202 1610 3224 1678
rect 3152 1594 3224 1610
rect 3254 1594 3304 1694
rect 3334 1678 3406 1694
rect 3334 1610 3356 1678
rect 3390 1610 3406 1678
rect 3334 1594 3406 1610
rect 3528 1678 3600 1694
rect 3528 1610 3544 1678
rect 3578 1610 3600 1678
rect 3528 1594 3600 1610
rect 3630 1678 3702 1694
rect 3630 1610 3652 1678
rect 3686 1610 3702 1678
rect 3630 1594 3702 1610
rect 3796 1678 3868 1694
rect 3796 1610 3812 1678
rect 3846 1610 3868 1678
rect 3796 1594 3868 1610
rect 3898 1594 3948 1694
rect 3978 1678 4050 1694
rect 3978 1610 4000 1678
rect 4034 1610 4050 1678
rect 3978 1594 4050 1610
rect 4132 1678 4204 1694
rect 4132 1610 4148 1678
rect 4182 1610 4204 1678
rect 4132 1594 4204 1610
rect 4234 1594 4284 1694
rect 4314 1678 4386 1694
rect 4314 1610 4336 1678
rect 4370 1610 4386 1678
rect 4314 1594 4386 1610
rect 4468 1678 4540 1694
rect 4468 1610 4484 1678
rect 4518 1610 4540 1678
rect 4468 1594 4540 1610
rect 4570 1678 4642 1694
rect 4570 1610 4592 1678
rect 4626 1610 4642 1678
rect 4570 1594 4642 1610
rect 4696 1678 4768 1694
rect 4696 1610 4712 1678
rect 4746 1610 4768 1678
rect 4696 1594 4768 1610
rect 4798 1594 4848 1694
rect 4878 1678 4950 1694
rect 4878 1610 4900 1678
rect 4934 1610 4950 1678
rect 4878 1594 4950 1610
rect 5032 1678 5104 1694
rect 5032 1610 5048 1678
rect 5082 1610 5104 1678
rect 5032 1594 5104 1610
rect 5134 1594 5184 1694
rect 5214 1678 5286 1694
rect 5214 1610 5236 1678
rect 5270 1610 5286 1678
rect 5214 1594 5286 1610
rect 5368 1678 5440 1694
rect 5368 1610 5384 1678
rect 5418 1610 5440 1678
rect 5368 1594 5440 1610
rect 5470 1594 5520 1694
rect 5550 1678 5622 1694
rect 5550 1610 5572 1678
rect 5606 1610 5622 1678
rect 5550 1594 5622 1610
rect 5704 1678 5776 1694
rect 5704 1610 5720 1678
rect 5754 1610 5776 1678
rect 5704 1594 5776 1610
rect 5806 1594 5856 1694
rect 5886 1678 5958 1694
rect 5886 1610 5908 1678
rect 5942 1610 5958 1678
rect 5886 1594 5958 1610
rect 6040 1678 6112 1694
rect 6040 1610 6056 1678
rect 6090 1610 6112 1678
rect 6040 1594 6112 1610
rect 6142 1678 6214 1694
rect 6142 1610 6164 1678
rect 6198 1610 6214 1678
rect 6142 1594 6214 1610
rect 6268 1678 6340 1694
rect 6268 1610 6284 1678
rect 6318 1610 6340 1678
rect 6268 1594 6340 1610
rect 6370 1594 6420 1694
rect 6450 1678 6522 1694
rect 6450 1610 6472 1678
rect 6506 1610 6522 1678
rect 6450 1594 6522 1610
rect 6604 1678 6676 1694
rect 6604 1610 6620 1678
rect 6654 1610 6676 1678
rect 6604 1594 6676 1610
rect 6706 1594 6756 1694
rect 6786 1678 6858 1694
rect 6786 1610 6808 1678
rect 6842 1610 6858 1678
rect 6786 1594 6858 1610
rect 6980 1678 7052 1694
rect 6980 1610 6996 1678
rect 7030 1610 7052 1678
rect 6980 1594 7052 1610
rect 7082 1678 7154 1694
rect 7082 1610 7104 1678
rect 7138 1610 7154 1678
rect 7082 1594 7154 1610
rect 7248 1678 7320 1694
rect 7248 1610 7264 1678
rect 7298 1610 7320 1678
rect 7248 1594 7320 1610
rect 7350 1594 7400 1694
rect 7430 1678 7502 1694
rect 7430 1610 7452 1678
rect 7486 1610 7502 1678
rect 7430 1594 7502 1610
rect 7584 1678 7656 1694
rect 7584 1610 7600 1678
rect 7634 1610 7656 1678
rect 7584 1594 7656 1610
rect 7686 1594 7736 1694
rect 7766 1678 7838 1694
rect 7766 1610 7788 1678
rect 7822 1610 7838 1678
rect 7766 1594 7838 1610
rect 7920 1678 7992 1694
rect 7920 1610 7936 1678
rect 7970 1610 7992 1678
rect 7920 1594 7992 1610
rect 8022 1678 8094 1694
rect 8022 1610 8044 1678
rect 8078 1610 8094 1678
rect 8022 1594 8094 1610
rect 8148 1678 8220 1694
rect 8148 1610 8164 1678
rect 8198 1610 8220 1678
rect 8148 1594 8220 1610
rect 8250 1594 8300 1694
rect 8330 1678 8402 1694
rect 8330 1610 8352 1678
rect 8386 1610 8402 1678
rect 8330 1594 8402 1610
rect 8484 1678 8556 1694
rect 8484 1610 8500 1678
rect 8534 1610 8556 1678
rect 8484 1594 8556 1610
rect 8586 1594 8636 1694
rect 8666 1678 8738 1694
rect 8666 1610 8688 1678
rect 8722 1610 8738 1678
rect 8666 1594 8738 1610
rect 8820 1678 8892 1694
rect 8820 1610 8836 1678
rect 8870 1610 8892 1678
rect 8820 1594 8892 1610
rect 8922 1594 8972 1694
rect 9002 1678 9074 1694
rect 9002 1610 9024 1678
rect 9058 1610 9074 1678
rect 9002 1594 9074 1610
rect 9156 1678 9228 1694
rect 9156 1610 9172 1678
rect 9206 1610 9228 1678
rect 9156 1594 9228 1610
rect 9258 1594 9308 1694
rect 9338 1678 9410 1694
rect 9338 1610 9360 1678
rect 9394 1610 9410 1678
rect 9338 1594 9410 1610
rect 9492 1678 9564 1694
rect 9492 1610 9508 1678
rect 9542 1610 9564 1678
rect 9492 1594 9564 1610
rect 9594 1678 9666 1694
rect 9594 1610 9616 1678
rect 9650 1610 9666 1678
rect 9594 1594 9666 1610
rect 9720 1678 9792 1694
rect 9720 1610 9736 1678
rect 9770 1610 9792 1678
rect 9720 1594 9792 1610
rect 9822 1594 9872 1694
rect 9902 1678 9974 1694
rect 9902 1610 9924 1678
rect 9958 1610 9974 1678
rect 9902 1594 9974 1610
rect 10056 1678 10128 1694
rect 10056 1610 10072 1678
rect 10106 1610 10128 1678
rect 10056 1594 10128 1610
rect 10158 1594 10208 1694
rect 10238 1678 10310 1694
rect 10238 1610 10260 1678
rect 10294 1610 10310 1678
rect 10238 1594 10310 1610
rect 10432 1678 10504 1694
rect 10432 1610 10448 1678
rect 10482 1610 10504 1678
rect 10432 1594 10504 1610
rect 10534 1678 10606 1694
rect 10534 1610 10556 1678
rect 10590 1610 10606 1678
rect 10534 1594 10606 1610
rect 10700 1678 10772 1694
rect 10700 1610 10716 1678
rect 10750 1610 10772 1678
rect 10700 1594 10772 1610
rect 10802 1594 10852 1694
rect 10882 1678 10954 1694
rect 10882 1610 10904 1678
rect 10938 1610 10954 1678
rect 10882 1594 10954 1610
rect 11036 1678 11108 1694
rect 11036 1610 11052 1678
rect 11086 1610 11108 1678
rect 11036 1594 11108 1610
rect 11138 1594 11188 1694
rect 11218 1678 11290 1694
rect 11218 1610 11240 1678
rect 11274 1610 11290 1678
rect 11218 1594 11290 1610
rect 11372 1678 11444 1694
rect 11372 1610 11388 1678
rect 11422 1610 11444 1678
rect 11372 1594 11444 1610
rect 11474 1678 11546 1694
rect 11474 1610 11496 1678
rect 11530 1610 11546 1678
rect 11474 1594 11546 1610
rect 11600 1678 11672 1694
rect 11600 1610 11616 1678
rect 11650 1610 11672 1678
rect 11600 1594 11672 1610
rect 11702 1594 11752 1694
rect 11782 1678 11854 1694
rect 11782 1610 11804 1678
rect 11838 1610 11854 1678
rect 11782 1594 11854 1610
rect 11936 1678 12008 1694
rect 11936 1610 11952 1678
rect 11986 1610 12008 1678
rect 11936 1594 12008 1610
rect 12038 1594 12088 1694
rect 12118 1678 12190 1694
rect 12118 1610 12140 1678
rect 12174 1610 12190 1678
rect 12118 1594 12190 1610
rect 12272 1678 12344 1694
rect 12272 1610 12288 1678
rect 12322 1610 12344 1678
rect 12272 1594 12344 1610
rect 12374 1594 12424 1694
rect 12454 1678 12526 1694
rect 12454 1610 12476 1678
rect 12510 1610 12526 1678
rect 12454 1594 12526 1610
rect 12608 1678 12680 1694
rect 12608 1610 12624 1678
rect 12658 1610 12680 1678
rect 12608 1594 12680 1610
rect 12710 1594 12760 1694
rect 12790 1678 12862 1694
rect 12790 1610 12812 1678
rect 12846 1610 12862 1678
rect 12790 1594 12862 1610
rect 12944 1678 13016 1694
rect 12944 1610 12960 1678
rect 12994 1610 13016 1678
rect 12944 1594 13016 1610
rect 13046 1678 13118 1694
rect 13046 1610 13068 1678
rect 13102 1610 13118 1678
rect 13046 1594 13118 1610
rect 13172 1678 13244 1694
rect 13172 1610 13188 1678
rect 13222 1610 13244 1678
rect 13172 1594 13244 1610
rect 13274 1594 13324 1694
rect 13354 1678 13426 1694
rect 13354 1610 13376 1678
rect 13410 1610 13426 1678
rect 13354 1594 13426 1610
rect 13508 1678 13580 1694
rect 13508 1610 13524 1678
rect 13558 1610 13580 1678
rect 13508 1594 13580 1610
rect 13610 1594 13660 1694
rect 13690 1678 13762 1694
rect 13690 1610 13712 1678
rect 13746 1610 13762 1678
rect 13690 1594 13762 1610
<< pdiff >>
rect 76 1178 148 1194
rect 76 1010 92 1178
rect 126 1010 148 1178
rect 76 994 148 1010
rect 178 1178 250 1194
rect 178 1010 200 1178
rect 234 1010 250 1178
rect 178 994 250 1010
rect 344 1178 416 1194
rect 344 1010 360 1178
rect 394 1010 416 1178
rect 344 994 416 1010
rect 446 1178 524 1194
rect 446 1010 468 1178
rect 502 1010 524 1178
rect 446 994 524 1010
rect 554 1178 626 1194
rect 554 1010 576 1178
rect 610 1010 626 1178
rect 554 994 626 1010
rect 680 1178 752 1194
rect 680 1010 696 1178
rect 730 1010 752 1178
rect 680 994 752 1010
rect 782 1178 860 1194
rect 782 1010 804 1178
rect 838 1010 860 1178
rect 782 994 860 1010
rect 890 1178 962 1194
rect 890 1010 912 1178
rect 946 1010 962 1178
rect 890 994 962 1010
rect 1016 1178 1088 1194
rect 1016 1010 1032 1178
rect 1066 1010 1088 1178
rect 1016 994 1088 1010
rect 1118 1178 1190 1194
rect 1118 1010 1140 1178
rect 1174 1010 1190 1178
rect 1118 994 1190 1010
rect 1244 1178 1316 1194
rect 1244 1010 1260 1178
rect 1294 1010 1316 1178
rect 1244 994 1316 1010
rect 1346 1178 1424 1194
rect 1346 1010 1368 1178
rect 1402 1010 1424 1178
rect 1346 994 1424 1010
rect 1454 1178 1526 1194
rect 1454 1010 1476 1178
rect 1510 1010 1526 1178
rect 1454 994 1526 1010
rect 1580 1178 1652 1194
rect 1580 1010 1596 1178
rect 1630 1010 1652 1178
rect 1580 994 1652 1010
rect 1682 1178 1760 1194
rect 1682 1010 1704 1178
rect 1738 1010 1760 1178
rect 1682 994 1760 1010
rect 1790 1178 1862 1194
rect 1790 1010 1812 1178
rect 1846 1010 1862 1178
rect 1790 994 1862 1010
rect 1916 1178 1988 1194
rect 1916 1010 1932 1178
rect 1966 1010 1988 1178
rect 1916 994 1988 1010
rect 2018 1178 2096 1194
rect 2018 1010 2040 1178
rect 2074 1010 2096 1178
rect 2018 994 2096 1010
rect 2126 1178 2198 1194
rect 2126 1010 2148 1178
rect 2182 1010 2198 1178
rect 2126 994 2198 1010
rect 2252 1178 2324 1194
rect 2252 1010 2268 1178
rect 2302 1010 2324 1178
rect 2252 994 2324 1010
rect 2354 1178 2432 1194
rect 2354 1010 2376 1178
rect 2410 1010 2432 1178
rect 2354 994 2432 1010
rect 2462 1178 2534 1194
rect 2462 1010 2484 1178
rect 2518 1010 2534 1178
rect 2462 994 2534 1010
rect 2588 1178 2660 1194
rect 2588 1010 2604 1178
rect 2638 1010 2660 1178
rect 2588 994 2660 1010
rect 2690 1178 2762 1194
rect 2690 1010 2712 1178
rect 2746 1010 2762 1178
rect 2690 994 2762 1010
rect 2816 1178 2888 1194
rect 2816 1010 2832 1178
rect 2866 1010 2888 1178
rect 2816 994 2888 1010
rect 2918 1178 2996 1194
rect 2918 1010 2940 1178
rect 2974 1010 2996 1178
rect 2918 994 2996 1010
rect 3026 1178 3098 1194
rect 3026 1010 3048 1178
rect 3082 1010 3098 1178
rect 3026 994 3098 1010
rect 3152 1178 3224 1194
rect 3152 1010 3168 1178
rect 3202 1010 3224 1178
rect 3152 994 3224 1010
rect 3254 1178 3332 1194
rect 3254 1010 3276 1178
rect 3310 1010 3332 1178
rect 3254 994 3332 1010
rect 3362 1178 3434 1194
rect 3362 1010 3384 1178
rect 3418 1010 3434 1178
rect 3362 994 3434 1010
rect 3528 1178 3600 1194
rect 3528 1010 3544 1178
rect 3578 1010 3600 1178
rect 3528 994 3600 1010
rect 3630 1178 3702 1194
rect 3630 1010 3652 1178
rect 3686 1010 3702 1178
rect 3630 994 3702 1010
rect 3796 1178 3868 1194
rect 3796 1010 3812 1178
rect 3846 1010 3868 1178
rect 3796 994 3868 1010
rect 3898 1178 3976 1194
rect 3898 1010 3920 1178
rect 3954 1010 3976 1178
rect 3898 994 3976 1010
rect 4006 1178 4078 1194
rect 4006 1010 4028 1178
rect 4062 1010 4078 1178
rect 4006 994 4078 1010
rect 4132 1178 4204 1194
rect 4132 1010 4148 1178
rect 4182 1010 4204 1178
rect 4132 994 4204 1010
rect 4234 1178 4312 1194
rect 4234 1010 4256 1178
rect 4290 1010 4312 1178
rect 4234 994 4312 1010
rect 4342 1178 4414 1194
rect 4342 1010 4364 1178
rect 4398 1010 4414 1178
rect 4342 994 4414 1010
rect 4468 1178 4540 1194
rect 4468 1010 4484 1178
rect 4518 1010 4540 1178
rect 4468 994 4540 1010
rect 4570 1178 4642 1194
rect 4570 1010 4592 1178
rect 4626 1010 4642 1178
rect 4570 994 4642 1010
rect 4696 1178 4768 1194
rect 4696 1010 4712 1178
rect 4746 1010 4768 1178
rect 4696 994 4768 1010
rect 4798 1178 4876 1194
rect 4798 1010 4820 1178
rect 4854 1010 4876 1178
rect 4798 994 4876 1010
rect 4906 1178 4978 1194
rect 4906 1010 4928 1178
rect 4962 1010 4978 1178
rect 4906 994 4978 1010
rect 5032 1178 5104 1194
rect 5032 1010 5048 1178
rect 5082 1010 5104 1178
rect 5032 994 5104 1010
rect 5134 1178 5212 1194
rect 5134 1010 5156 1178
rect 5190 1010 5212 1178
rect 5134 994 5212 1010
rect 5242 1178 5314 1194
rect 5242 1010 5264 1178
rect 5298 1010 5314 1178
rect 5242 994 5314 1010
rect 5368 1178 5440 1194
rect 5368 1010 5384 1178
rect 5418 1010 5440 1178
rect 5368 994 5440 1010
rect 5470 1178 5548 1194
rect 5470 1010 5492 1178
rect 5526 1010 5548 1178
rect 5470 994 5548 1010
rect 5578 1178 5650 1194
rect 5578 1010 5600 1178
rect 5634 1010 5650 1178
rect 5578 994 5650 1010
rect 5704 1178 5776 1194
rect 5704 1010 5720 1178
rect 5754 1010 5776 1178
rect 5704 994 5776 1010
rect 5806 1178 5884 1194
rect 5806 1010 5828 1178
rect 5862 1010 5884 1178
rect 5806 994 5884 1010
rect 5914 1178 5986 1194
rect 5914 1010 5936 1178
rect 5970 1010 5986 1178
rect 5914 994 5986 1010
rect 6040 1178 6112 1194
rect 6040 1010 6056 1178
rect 6090 1010 6112 1178
rect 6040 994 6112 1010
rect 6142 1178 6214 1194
rect 6142 1010 6164 1178
rect 6198 1010 6214 1178
rect 6142 994 6214 1010
rect 6268 1178 6340 1194
rect 6268 1010 6284 1178
rect 6318 1010 6340 1178
rect 6268 994 6340 1010
rect 6370 1178 6448 1194
rect 6370 1010 6392 1178
rect 6426 1010 6448 1178
rect 6370 994 6448 1010
rect 6478 1178 6550 1194
rect 6478 1010 6500 1178
rect 6534 1010 6550 1178
rect 6478 994 6550 1010
rect 6604 1178 6676 1194
rect 6604 1010 6620 1178
rect 6654 1010 6676 1178
rect 6604 994 6676 1010
rect 6706 1178 6784 1194
rect 6706 1010 6728 1178
rect 6762 1010 6784 1178
rect 6706 994 6784 1010
rect 6814 1178 6886 1194
rect 6814 1010 6836 1178
rect 6870 1010 6886 1178
rect 6814 994 6886 1010
rect 6980 1178 7052 1194
rect 6980 1010 6996 1178
rect 7030 1010 7052 1178
rect 6980 994 7052 1010
rect 7082 1178 7154 1194
rect 7082 1010 7104 1178
rect 7138 1010 7154 1178
rect 7082 994 7154 1010
rect 7248 1178 7320 1194
rect 7248 1010 7264 1178
rect 7298 1010 7320 1178
rect 7248 994 7320 1010
rect 7350 1178 7428 1194
rect 7350 1010 7372 1178
rect 7406 1010 7428 1178
rect 7350 994 7428 1010
rect 7458 1178 7530 1194
rect 7458 1010 7480 1178
rect 7514 1010 7530 1178
rect 7458 994 7530 1010
rect 7584 1178 7656 1194
rect 7584 1010 7600 1178
rect 7634 1010 7656 1178
rect 7584 994 7656 1010
rect 7686 1178 7764 1194
rect 7686 1010 7708 1178
rect 7742 1010 7764 1178
rect 7686 994 7764 1010
rect 7794 1178 7866 1194
rect 7794 1010 7816 1178
rect 7850 1010 7866 1178
rect 7794 994 7866 1010
rect 7920 1178 7992 1194
rect 7920 1010 7936 1178
rect 7970 1010 7992 1178
rect 7920 994 7992 1010
rect 8022 1178 8094 1194
rect 8022 1010 8044 1178
rect 8078 1010 8094 1178
rect 8022 994 8094 1010
rect 8148 1178 8220 1194
rect 8148 1010 8164 1178
rect 8198 1010 8220 1178
rect 8148 994 8220 1010
rect 8250 1178 8328 1194
rect 8250 1010 8272 1178
rect 8306 1010 8328 1178
rect 8250 994 8328 1010
rect 8358 1178 8430 1194
rect 8358 1010 8380 1178
rect 8414 1010 8430 1178
rect 8358 994 8430 1010
rect 8484 1178 8556 1194
rect 8484 1010 8500 1178
rect 8534 1010 8556 1178
rect 8484 994 8556 1010
rect 8586 1178 8664 1194
rect 8586 1010 8608 1178
rect 8642 1010 8664 1178
rect 8586 994 8664 1010
rect 8694 1178 8766 1194
rect 8694 1010 8716 1178
rect 8750 1010 8766 1178
rect 8694 994 8766 1010
rect 8820 1178 8892 1194
rect 8820 1010 8836 1178
rect 8870 1010 8892 1178
rect 8820 994 8892 1010
rect 8922 1178 9000 1194
rect 8922 1010 8944 1178
rect 8978 1010 9000 1178
rect 8922 994 9000 1010
rect 9030 1178 9102 1194
rect 9030 1010 9052 1178
rect 9086 1010 9102 1178
rect 9030 994 9102 1010
rect 9156 1178 9228 1194
rect 9156 1010 9172 1178
rect 9206 1010 9228 1178
rect 9156 994 9228 1010
rect 9258 1178 9336 1194
rect 9258 1010 9280 1178
rect 9314 1010 9336 1178
rect 9258 994 9336 1010
rect 9366 1178 9438 1194
rect 9366 1010 9388 1178
rect 9422 1010 9438 1178
rect 9366 994 9438 1010
rect 9492 1178 9564 1194
rect 9492 1010 9508 1178
rect 9542 1010 9564 1178
rect 9492 994 9564 1010
rect 9594 1178 9666 1194
rect 9594 1010 9616 1178
rect 9650 1010 9666 1178
rect 9594 994 9666 1010
rect 9720 1178 9792 1194
rect 9720 1010 9736 1178
rect 9770 1010 9792 1178
rect 9720 994 9792 1010
rect 9822 1178 9900 1194
rect 9822 1010 9844 1178
rect 9878 1010 9900 1178
rect 9822 994 9900 1010
rect 9930 1178 10002 1194
rect 9930 1010 9952 1178
rect 9986 1010 10002 1178
rect 9930 994 10002 1010
rect 10056 1178 10128 1194
rect 10056 1010 10072 1178
rect 10106 1010 10128 1178
rect 10056 994 10128 1010
rect 10158 1178 10236 1194
rect 10158 1010 10180 1178
rect 10214 1010 10236 1178
rect 10158 994 10236 1010
rect 10266 1178 10338 1194
rect 10266 1010 10288 1178
rect 10322 1010 10338 1178
rect 10266 994 10338 1010
rect 10432 1178 10504 1194
rect 10432 1010 10448 1178
rect 10482 1010 10504 1178
rect 10432 994 10504 1010
rect 10534 1178 10606 1194
rect 10534 1010 10556 1178
rect 10590 1010 10606 1178
rect 10534 994 10606 1010
rect 10700 1178 10772 1194
rect 10700 1010 10716 1178
rect 10750 1010 10772 1178
rect 10700 994 10772 1010
rect 10802 1178 10880 1194
rect 10802 1010 10824 1178
rect 10858 1010 10880 1178
rect 10802 994 10880 1010
rect 10910 1178 10982 1194
rect 10910 1010 10932 1178
rect 10966 1010 10982 1178
rect 10910 994 10982 1010
rect 11036 1178 11108 1194
rect 11036 1010 11052 1178
rect 11086 1010 11108 1178
rect 11036 994 11108 1010
rect 11138 1178 11216 1194
rect 11138 1010 11160 1178
rect 11194 1010 11216 1178
rect 11138 994 11216 1010
rect 11246 1178 11318 1194
rect 11246 1010 11268 1178
rect 11302 1010 11318 1178
rect 11246 994 11318 1010
rect 11372 1178 11444 1194
rect 11372 1010 11388 1178
rect 11422 1010 11444 1178
rect 11372 994 11444 1010
rect 11474 1178 11546 1194
rect 11474 1010 11496 1178
rect 11530 1010 11546 1178
rect 11474 994 11546 1010
rect 11600 1178 11672 1194
rect 11600 1010 11616 1178
rect 11650 1010 11672 1178
rect 11600 994 11672 1010
rect 11702 1178 11780 1194
rect 11702 1010 11724 1178
rect 11758 1010 11780 1178
rect 11702 994 11780 1010
rect 11810 1178 11882 1194
rect 11810 1010 11832 1178
rect 11866 1010 11882 1178
rect 11810 994 11882 1010
rect 11936 1178 12008 1194
rect 11936 1010 11952 1178
rect 11986 1010 12008 1178
rect 11936 994 12008 1010
rect 12038 1178 12116 1194
rect 12038 1010 12060 1178
rect 12094 1010 12116 1178
rect 12038 994 12116 1010
rect 12146 1178 12218 1194
rect 12146 1010 12168 1178
rect 12202 1010 12218 1178
rect 12146 994 12218 1010
rect 12272 1178 12344 1194
rect 12272 1010 12288 1178
rect 12322 1010 12344 1178
rect 12272 994 12344 1010
rect 12374 1178 12452 1194
rect 12374 1010 12396 1178
rect 12430 1010 12452 1178
rect 12374 994 12452 1010
rect 12482 1178 12554 1194
rect 12482 1010 12504 1178
rect 12538 1010 12554 1178
rect 12482 994 12554 1010
rect 12608 1178 12680 1194
rect 12608 1010 12624 1178
rect 12658 1010 12680 1178
rect 12608 994 12680 1010
rect 12710 1178 12788 1194
rect 12710 1010 12732 1178
rect 12766 1010 12788 1178
rect 12710 994 12788 1010
rect 12818 1178 12890 1194
rect 12818 1010 12840 1178
rect 12874 1010 12890 1178
rect 12818 994 12890 1010
rect 12944 1178 13016 1194
rect 12944 1010 12960 1178
rect 12994 1010 13016 1178
rect 12944 994 13016 1010
rect 13046 1178 13118 1194
rect 13046 1010 13068 1178
rect 13102 1010 13118 1178
rect 13046 994 13118 1010
rect 13172 1178 13244 1194
rect 13172 1010 13188 1178
rect 13222 1010 13244 1178
rect 13172 994 13244 1010
rect 13274 1178 13352 1194
rect 13274 1010 13296 1178
rect 13330 1010 13352 1178
rect 13274 994 13352 1010
rect 13382 1178 13454 1194
rect 13382 1010 13404 1178
rect 13438 1010 13454 1178
rect 13382 994 13454 1010
rect 13508 1178 13580 1194
rect 13508 1010 13524 1178
rect 13558 1010 13580 1178
rect 13508 994 13580 1010
rect 13610 1178 13688 1194
rect 13610 1010 13632 1178
rect 13666 1010 13688 1178
rect 13610 994 13688 1010
rect 13718 1178 13790 1194
rect 13718 1010 13740 1178
rect 13774 1010 13790 1178
rect 13718 994 13790 1010
<< ndiffc >>
rect 92 1610 126 1678
rect 200 1610 234 1678
rect 360 1610 394 1678
rect 548 1610 582 1678
rect 696 1610 730 1678
rect 884 1610 918 1678
rect 1032 1610 1066 1678
rect 1140 1610 1174 1678
rect 1260 1610 1294 1678
rect 1448 1610 1482 1678
rect 1596 1610 1630 1678
rect 1784 1610 1818 1678
rect 1932 1610 1966 1678
rect 2120 1610 2154 1678
rect 2268 1610 2302 1678
rect 2456 1610 2490 1678
rect 2604 1610 2638 1678
rect 2712 1610 2746 1678
rect 2832 1610 2866 1678
rect 3020 1610 3054 1678
rect 3168 1610 3202 1678
rect 3356 1610 3390 1678
rect 3544 1610 3578 1678
rect 3652 1610 3686 1678
rect 3812 1610 3846 1678
rect 4000 1610 4034 1678
rect 4148 1610 4182 1678
rect 4336 1610 4370 1678
rect 4484 1610 4518 1678
rect 4592 1610 4626 1678
rect 4712 1610 4746 1678
rect 4900 1610 4934 1678
rect 5048 1610 5082 1678
rect 5236 1610 5270 1678
rect 5384 1610 5418 1678
rect 5572 1610 5606 1678
rect 5720 1610 5754 1678
rect 5908 1610 5942 1678
rect 6056 1610 6090 1678
rect 6164 1610 6198 1678
rect 6284 1610 6318 1678
rect 6472 1610 6506 1678
rect 6620 1610 6654 1678
rect 6808 1610 6842 1678
rect 6996 1610 7030 1678
rect 7104 1610 7138 1678
rect 7264 1610 7298 1678
rect 7452 1610 7486 1678
rect 7600 1610 7634 1678
rect 7788 1610 7822 1678
rect 7936 1610 7970 1678
rect 8044 1610 8078 1678
rect 8164 1610 8198 1678
rect 8352 1610 8386 1678
rect 8500 1610 8534 1678
rect 8688 1610 8722 1678
rect 8836 1610 8870 1678
rect 9024 1610 9058 1678
rect 9172 1610 9206 1678
rect 9360 1610 9394 1678
rect 9508 1610 9542 1678
rect 9616 1610 9650 1678
rect 9736 1610 9770 1678
rect 9924 1610 9958 1678
rect 10072 1610 10106 1678
rect 10260 1610 10294 1678
rect 10448 1610 10482 1678
rect 10556 1610 10590 1678
rect 10716 1610 10750 1678
rect 10904 1610 10938 1678
rect 11052 1610 11086 1678
rect 11240 1610 11274 1678
rect 11388 1610 11422 1678
rect 11496 1610 11530 1678
rect 11616 1610 11650 1678
rect 11804 1610 11838 1678
rect 11952 1610 11986 1678
rect 12140 1610 12174 1678
rect 12288 1610 12322 1678
rect 12476 1610 12510 1678
rect 12624 1610 12658 1678
rect 12812 1610 12846 1678
rect 12960 1610 12994 1678
rect 13068 1610 13102 1678
rect 13188 1610 13222 1678
rect 13376 1610 13410 1678
rect 13524 1610 13558 1678
rect 13712 1610 13746 1678
<< pdiffc >>
rect 92 1010 126 1178
rect 200 1010 234 1178
rect 360 1010 394 1178
rect 468 1010 502 1178
rect 576 1010 610 1178
rect 696 1010 730 1178
rect 804 1010 838 1178
rect 912 1010 946 1178
rect 1032 1010 1066 1178
rect 1140 1010 1174 1178
rect 1260 1010 1294 1178
rect 1368 1010 1402 1178
rect 1476 1010 1510 1178
rect 1596 1010 1630 1178
rect 1704 1010 1738 1178
rect 1812 1010 1846 1178
rect 1932 1010 1966 1178
rect 2040 1010 2074 1178
rect 2148 1010 2182 1178
rect 2268 1010 2302 1178
rect 2376 1010 2410 1178
rect 2484 1010 2518 1178
rect 2604 1010 2638 1178
rect 2712 1010 2746 1178
rect 2832 1010 2866 1178
rect 2940 1010 2974 1178
rect 3048 1010 3082 1178
rect 3168 1010 3202 1178
rect 3276 1010 3310 1178
rect 3384 1010 3418 1178
rect 3544 1010 3578 1178
rect 3652 1010 3686 1178
rect 3812 1010 3846 1178
rect 3920 1010 3954 1178
rect 4028 1010 4062 1178
rect 4148 1010 4182 1178
rect 4256 1010 4290 1178
rect 4364 1010 4398 1178
rect 4484 1010 4518 1178
rect 4592 1010 4626 1178
rect 4712 1010 4746 1178
rect 4820 1010 4854 1178
rect 4928 1010 4962 1178
rect 5048 1010 5082 1178
rect 5156 1010 5190 1178
rect 5264 1010 5298 1178
rect 5384 1010 5418 1178
rect 5492 1010 5526 1178
rect 5600 1010 5634 1178
rect 5720 1010 5754 1178
rect 5828 1010 5862 1178
rect 5936 1010 5970 1178
rect 6056 1010 6090 1178
rect 6164 1010 6198 1178
rect 6284 1010 6318 1178
rect 6392 1010 6426 1178
rect 6500 1010 6534 1178
rect 6620 1010 6654 1178
rect 6728 1010 6762 1178
rect 6836 1010 6870 1178
rect 6996 1010 7030 1178
rect 7104 1010 7138 1178
rect 7264 1010 7298 1178
rect 7372 1010 7406 1178
rect 7480 1010 7514 1178
rect 7600 1010 7634 1178
rect 7708 1010 7742 1178
rect 7816 1010 7850 1178
rect 7936 1010 7970 1178
rect 8044 1010 8078 1178
rect 8164 1010 8198 1178
rect 8272 1010 8306 1178
rect 8380 1010 8414 1178
rect 8500 1010 8534 1178
rect 8608 1010 8642 1178
rect 8716 1010 8750 1178
rect 8836 1010 8870 1178
rect 8944 1010 8978 1178
rect 9052 1010 9086 1178
rect 9172 1010 9206 1178
rect 9280 1010 9314 1178
rect 9388 1010 9422 1178
rect 9508 1010 9542 1178
rect 9616 1010 9650 1178
rect 9736 1010 9770 1178
rect 9844 1010 9878 1178
rect 9952 1010 9986 1178
rect 10072 1010 10106 1178
rect 10180 1010 10214 1178
rect 10288 1010 10322 1178
rect 10448 1010 10482 1178
rect 10556 1010 10590 1178
rect 10716 1010 10750 1178
rect 10824 1010 10858 1178
rect 10932 1010 10966 1178
rect 11052 1010 11086 1178
rect 11160 1010 11194 1178
rect 11268 1010 11302 1178
rect 11388 1010 11422 1178
rect 11496 1010 11530 1178
rect 11616 1010 11650 1178
rect 11724 1010 11758 1178
rect 11832 1010 11866 1178
rect 11952 1010 11986 1178
rect 12060 1010 12094 1178
rect 12168 1010 12202 1178
rect 12288 1010 12322 1178
rect 12396 1010 12430 1178
rect 12504 1010 12538 1178
rect 12624 1010 12658 1178
rect 12732 1010 12766 1178
rect 12840 1010 12874 1178
rect 12960 1010 12994 1178
rect 13068 1010 13102 1178
rect 13188 1010 13222 1178
rect 13296 1010 13330 1178
rect 13404 1010 13438 1178
rect 13524 1010 13558 1178
rect 13632 1010 13666 1178
rect 13740 1010 13774 1178
<< psubdiff >>
rect 36 1748 60 1804
rect 266 1748 290 1804
rect 344 1748 368 1804
rect 1810 1748 1834 1804
rect 1916 1748 1940 1804
rect 3382 1748 3406 1804
rect 3488 1748 3512 1804
rect 3718 1748 3742 1804
rect 3796 1748 3820 1804
rect 5262 1748 5286 1804
rect 5368 1748 5392 1804
rect 6834 1748 6858 1804
rect 6940 1748 6964 1804
rect 7170 1748 7194 1804
rect 7248 1748 7272 1804
rect 8714 1748 8738 1804
rect 8820 1748 8844 1804
rect 10286 1748 10310 1804
rect 10392 1748 10416 1804
rect 10622 1748 10646 1804
rect 10700 1748 10724 1804
rect 12166 1748 12190 1804
rect 12272 1748 12296 1804
rect 13738 1748 13762 1804
<< nsubdiff >>
rect 36 884 60 940
rect 266 884 290 940
rect 344 884 368 940
rect 1838 884 1862 940
rect 1916 884 1940 940
rect 3410 884 3434 940
rect 3488 884 3512 940
rect 3718 884 3742 940
rect 3796 884 3820 940
rect 5290 884 5314 940
rect 5368 884 5392 940
rect 6862 884 6886 940
rect 6940 884 6964 940
rect 7170 884 7194 940
rect 7248 884 7272 940
rect 8742 884 8766 940
rect 8820 884 8844 940
rect 10314 884 10338 940
rect 10392 884 10416 940
rect 10622 884 10646 940
rect 10700 884 10724 940
rect 12194 884 12218 940
rect 12272 884 12296 940
rect 13766 884 13790 940
<< psubdiffcont >>
rect 60 1748 266 1804
rect 368 1748 1810 1804
rect 1940 1748 3382 1804
rect 3512 1748 3718 1804
rect 3820 1748 5262 1804
rect 5392 1748 6834 1804
rect 6964 1748 7170 1804
rect 7272 1748 8714 1804
rect 8844 1748 10286 1804
rect 10416 1748 10622 1804
rect 10724 1748 12166 1804
rect 12296 1748 13738 1804
<< nsubdiffcont >>
rect 60 884 266 940
rect 368 884 1838 940
rect 1940 884 3410 940
rect 3512 884 3718 940
rect 3820 884 5290 940
rect 5392 884 6862 940
rect 6964 884 7170 940
rect 7272 884 8742 940
rect 8844 884 10314 940
rect 10416 884 10622 940
rect 10724 884 12194 940
rect 12296 884 13766 940
<< poly >>
rect 148 1694 178 1720
rect 416 1694 446 1720
rect 496 1694 526 1720
rect 752 1694 782 1720
rect 832 1694 862 1720
rect 1088 1694 1118 1720
rect 1316 1694 1346 1720
rect 1396 1694 1426 1720
rect 1652 1694 1682 1720
rect 1732 1694 1762 1720
rect 1988 1694 2018 1720
rect 2068 1694 2098 1720
rect 2324 1694 2354 1720
rect 2404 1694 2434 1720
rect 2660 1694 2690 1720
rect 2888 1694 2918 1720
rect 2968 1694 2998 1720
rect 3224 1694 3254 1720
rect 3304 1694 3334 1720
rect 3600 1694 3630 1720
rect 3868 1694 3898 1720
rect 3948 1694 3978 1720
rect 4204 1694 4234 1720
rect 4284 1694 4314 1720
rect 4540 1694 4570 1720
rect 4768 1694 4798 1720
rect 4848 1694 4878 1720
rect 5104 1694 5134 1720
rect 5184 1694 5214 1720
rect 5440 1694 5470 1720
rect 5520 1694 5550 1720
rect 5776 1694 5806 1720
rect 5856 1694 5886 1720
rect 6112 1694 6142 1720
rect 6340 1694 6370 1720
rect 6420 1694 6450 1720
rect 6676 1694 6706 1720
rect 6756 1694 6786 1720
rect 7052 1694 7082 1720
rect 7320 1694 7350 1720
rect 7400 1694 7430 1720
rect 7656 1694 7686 1720
rect 7736 1694 7766 1720
rect 7992 1694 8022 1720
rect 8220 1694 8250 1720
rect 8300 1694 8330 1720
rect 8556 1694 8586 1720
rect 8636 1694 8666 1720
rect 8892 1694 8922 1720
rect 8972 1694 9002 1720
rect 9228 1694 9258 1720
rect 9308 1694 9338 1720
rect 9564 1694 9594 1720
rect 9792 1694 9822 1720
rect 9872 1694 9902 1720
rect 10128 1694 10158 1720
rect 10208 1694 10238 1720
rect 10504 1694 10534 1720
rect 10772 1694 10802 1720
rect 10852 1694 10882 1720
rect 11108 1694 11138 1720
rect 11188 1694 11218 1720
rect 11444 1694 11474 1720
rect 11672 1694 11702 1720
rect 11752 1694 11782 1720
rect 12008 1694 12038 1720
rect 12088 1694 12118 1720
rect 12344 1694 12374 1720
rect 12424 1694 12454 1720
rect 12680 1694 12710 1720
rect 12760 1694 12790 1720
rect 13016 1694 13046 1720
rect 13244 1694 13274 1720
rect 13324 1694 13354 1720
rect 13580 1694 13610 1720
rect 13660 1694 13690 1720
rect 148 1426 178 1594
rect 82 1410 178 1426
rect 82 1376 98 1410
rect 132 1376 178 1410
rect 82 1360 178 1376
rect 148 1194 178 1360
rect 416 1296 446 1594
rect 496 1532 526 1594
rect 496 1502 554 1532
rect 350 1280 446 1296
rect 350 1246 366 1280
rect 400 1246 446 1280
rect 350 1230 446 1246
rect 416 1194 446 1230
rect 524 1396 554 1502
rect 752 1396 782 1594
rect 832 1532 862 1594
rect 832 1502 890 1532
rect 524 1380 782 1396
rect 524 1346 634 1380
rect 668 1346 782 1380
rect 524 1330 782 1346
rect 524 1194 554 1330
rect 752 1194 782 1330
rect 860 1396 890 1502
rect 860 1380 956 1396
rect 860 1346 906 1380
rect 940 1346 956 1380
rect 860 1330 956 1346
rect 860 1194 890 1330
rect 1088 1296 1118 1594
rect 1316 1426 1346 1594
rect 1396 1532 1426 1594
rect 1396 1502 1454 1532
rect 1250 1410 1346 1426
rect 1250 1376 1266 1410
rect 1300 1376 1346 1410
rect 1250 1360 1346 1376
rect 1022 1280 1118 1296
rect 1022 1246 1038 1280
rect 1072 1246 1118 1280
rect 1022 1230 1118 1246
rect 1088 1194 1118 1230
rect 1316 1194 1346 1360
rect 1424 1344 1454 1502
rect 1652 1426 1682 1594
rect 1732 1532 1762 1594
rect 1732 1502 1790 1532
rect 1586 1410 1682 1426
rect 1586 1376 1602 1410
rect 1636 1376 1682 1410
rect 1586 1360 1682 1376
rect 1424 1328 1520 1344
rect 1424 1294 1470 1328
rect 1504 1294 1520 1328
rect 1424 1278 1520 1294
rect 1424 1194 1454 1278
rect 1652 1194 1682 1360
rect 1760 1344 1790 1502
rect 1760 1328 1856 1344
rect 1760 1294 1806 1328
rect 1840 1294 1856 1328
rect 1988 1296 2018 1594
rect 2068 1532 2098 1594
rect 2068 1502 2126 1532
rect 1760 1278 1856 1294
rect 1922 1280 2018 1296
rect 1760 1194 1790 1278
rect 1922 1246 1938 1280
rect 1972 1246 2018 1280
rect 1922 1230 2018 1246
rect 1988 1194 2018 1230
rect 2096 1396 2126 1502
rect 2324 1396 2354 1594
rect 2404 1532 2434 1594
rect 2404 1502 2462 1532
rect 2096 1380 2354 1396
rect 2096 1346 2206 1380
rect 2240 1346 2354 1380
rect 2096 1330 2354 1346
rect 2096 1194 2126 1330
rect 2324 1194 2354 1330
rect 2432 1396 2462 1502
rect 2432 1380 2528 1396
rect 2432 1346 2478 1380
rect 2512 1346 2528 1380
rect 2432 1330 2528 1346
rect 2432 1194 2462 1330
rect 2660 1296 2690 1594
rect 2888 1426 2918 1594
rect 2968 1532 2998 1594
rect 2968 1502 3026 1532
rect 2822 1410 2918 1426
rect 2822 1376 2838 1410
rect 2872 1376 2918 1410
rect 2822 1360 2918 1376
rect 2594 1280 2690 1296
rect 2594 1246 2610 1280
rect 2644 1246 2690 1280
rect 2594 1230 2690 1246
rect 2660 1194 2690 1230
rect 2888 1194 2918 1360
rect 2996 1344 3026 1502
rect 3224 1426 3254 1594
rect 3304 1532 3334 1594
rect 3304 1502 3362 1532
rect 3158 1410 3254 1426
rect 3158 1376 3174 1410
rect 3208 1376 3254 1410
rect 3158 1360 3254 1376
rect 2996 1328 3092 1344
rect 2996 1294 3042 1328
rect 3076 1294 3092 1328
rect 2996 1278 3092 1294
rect 2996 1194 3026 1278
rect 3224 1194 3254 1360
rect 3332 1344 3362 1502
rect 3600 1426 3630 1594
rect 3534 1410 3630 1426
rect 3534 1376 3550 1410
rect 3584 1376 3630 1410
rect 3534 1360 3630 1376
rect 3332 1328 3428 1344
rect 3332 1294 3378 1328
rect 3412 1294 3428 1328
rect 3332 1278 3428 1294
rect 3332 1194 3362 1278
rect 3600 1194 3630 1360
rect 3868 1296 3898 1594
rect 3948 1532 3978 1594
rect 3948 1502 4006 1532
rect 3802 1280 3898 1296
rect 3802 1246 3818 1280
rect 3852 1246 3898 1280
rect 3802 1230 3898 1246
rect 3868 1194 3898 1230
rect 3976 1396 4006 1502
rect 4204 1396 4234 1594
rect 4284 1532 4314 1594
rect 4284 1502 4342 1532
rect 3976 1380 4234 1396
rect 3976 1346 4086 1380
rect 4120 1346 4234 1380
rect 3976 1330 4234 1346
rect 3976 1194 4006 1330
rect 4204 1194 4234 1330
rect 4312 1396 4342 1502
rect 4312 1380 4408 1396
rect 4312 1346 4358 1380
rect 4392 1346 4408 1380
rect 4312 1330 4408 1346
rect 4312 1194 4342 1330
rect 4540 1296 4570 1594
rect 4768 1426 4798 1594
rect 4848 1532 4878 1594
rect 4848 1502 4906 1532
rect 4702 1410 4798 1426
rect 4702 1376 4718 1410
rect 4752 1376 4798 1410
rect 4702 1360 4798 1376
rect 4474 1280 4570 1296
rect 4474 1246 4490 1280
rect 4524 1246 4570 1280
rect 4474 1230 4570 1246
rect 4540 1194 4570 1230
rect 4768 1194 4798 1360
rect 4876 1344 4906 1502
rect 5104 1426 5134 1594
rect 5184 1532 5214 1594
rect 5184 1502 5242 1532
rect 5038 1410 5134 1426
rect 5038 1376 5054 1410
rect 5088 1376 5134 1410
rect 5038 1360 5134 1376
rect 4876 1328 4972 1344
rect 4876 1294 4922 1328
rect 4956 1294 4972 1328
rect 4876 1278 4972 1294
rect 4876 1194 4906 1278
rect 5104 1194 5134 1360
rect 5212 1344 5242 1502
rect 5212 1328 5308 1344
rect 5212 1294 5258 1328
rect 5292 1294 5308 1328
rect 5440 1296 5470 1594
rect 5520 1532 5550 1594
rect 5520 1502 5578 1532
rect 5212 1278 5308 1294
rect 5374 1280 5470 1296
rect 5212 1194 5242 1278
rect 5374 1246 5390 1280
rect 5424 1246 5470 1280
rect 5374 1230 5470 1246
rect 5440 1194 5470 1230
rect 5548 1396 5578 1502
rect 5776 1396 5806 1594
rect 5856 1532 5886 1594
rect 5856 1502 5914 1532
rect 5548 1380 5806 1396
rect 5548 1346 5658 1380
rect 5692 1346 5806 1380
rect 5548 1330 5806 1346
rect 5548 1194 5578 1330
rect 5776 1194 5806 1330
rect 5884 1396 5914 1502
rect 5884 1380 5980 1396
rect 5884 1346 5930 1380
rect 5964 1346 5980 1380
rect 5884 1330 5980 1346
rect 5884 1194 5914 1330
rect 6112 1296 6142 1594
rect 6340 1426 6370 1594
rect 6420 1532 6450 1594
rect 6420 1502 6478 1532
rect 6274 1410 6370 1426
rect 6274 1376 6290 1410
rect 6324 1376 6370 1410
rect 6274 1360 6370 1376
rect 6046 1280 6142 1296
rect 6046 1246 6062 1280
rect 6096 1246 6142 1280
rect 6046 1230 6142 1246
rect 6112 1194 6142 1230
rect 6340 1194 6370 1360
rect 6448 1344 6478 1502
rect 6676 1426 6706 1594
rect 6756 1532 6786 1594
rect 6756 1502 6814 1532
rect 6610 1410 6706 1426
rect 6610 1376 6626 1410
rect 6660 1376 6706 1410
rect 6610 1360 6706 1376
rect 6448 1328 6544 1344
rect 6448 1294 6494 1328
rect 6528 1294 6544 1328
rect 6448 1278 6544 1294
rect 6448 1194 6478 1278
rect 6676 1194 6706 1360
rect 6784 1344 6814 1502
rect 7052 1426 7082 1594
rect 6986 1410 7082 1426
rect 6986 1376 7002 1410
rect 7036 1376 7082 1410
rect 6986 1360 7082 1376
rect 6784 1328 6880 1344
rect 6784 1294 6830 1328
rect 6864 1294 6880 1328
rect 6784 1278 6880 1294
rect 6784 1194 6814 1278
rect 7052 1194 7082 1360
rect 7320 1296 7350 1594
rect 7400 1532 7430 1594
rect 7400 1502 7458 1532
rect 7254 1280 7350 1296
rect 7254 1246 7270 1280
rect 7304 1246 7350 1280
rect 7254 1230 7350 1246
rect 7320 1194 7350 1230
rect 7428 1396 7458 1502
rect 7656 1396 7686 1594
rect 7736 1532 7766 1594
rect 7736 1502 7794 1532
rect 7428 1380 7686 1396
rect 7428 1346 7538 1380
rect 7572 1346 7686 1380
rect 7428 1330 7686 1346
rect 7428 1194 7458 1330
rect 7656 1194 7686 1330
rect 7764 1396 7794 1502
rect 7764 1380 7860 1396
rect 7764 1346 7810 1380
rect 7844 1346 7860 1380
rect 7764 1330 7860 1346
rect 7764 1194 7794 1330
rect 7992 1296 8022 1594
rect 8220 1426 8250 1594
rect 8300 1532 8330 1594
rect 8300 1502 8358 1532
rect 8154 1410 8250 1426
rect 8154 1376 8170 1410
rect 8204 1376 8250 1410
rect 8154 1360 8250 1376
rect 7926 1280 8022 1296
rect 7926 1246 7942 1280
rect 7976 1246 8022 1280
rect 7926 1230 8022 1246
rect 7992 1194 8022 1230
rect 8220 1194 8250 1360
rect 8328 1344 8358 1502
rect 8556 1426 8586 1594
rect 8636 1532 8666 1594
rect 8636 1502 8694 1532
rect 8490 1410 8586 1426
rect 8490 1376 8506 1410
rect 8540 1376 8586 1410
rect 8490 1360 8586 1376
rect 8328 1328 8424 1344
rect 8328 1294 8374 1328
rect 8408 1294 8424 1328
rect 8328 1278 8424 1294
rect 8328 1194 8358 1278
rect 8556 1194 8586 1360
rect 8664 1344 8694 1502
rect 8664 1328 8760 1344
rect 8664 1294 8710 1328
rect 8744 1294 8760 1328
rect 8892 1296 8922 1594
rect 8972 1532 9002 1594
rect 8972 1502 9030 1532
rect 8664 1278 8760 1294
rect 8826 1280 8922 1296
rect 8664 1194 8694 1278
rect 8826 1246 8842 1280
rect 8876 1246 8922 1280
rect 8826 1230 8922 1246
rect 8892 1194 8922 1230
rect 9000 1396 9030 1502
rect 9228 1396 9258 1594
rect 9308 1532 9338 1594
rect 9308 1502 9366 1532
rect 9000 1380 9258 1396
rect 9000 1346 9110 1380
rect 9144 1346 9258 1380
rect 9000 1330 9258 1346
rect 9000 1194 9030 1330
rect 9228 1194 9258 1330
rect 9336 1396 9366 1502
rect 9336 1380 9432 1396
rect 9336 1346 9382 1380
rect 9416 1346 9432 1380
rect 9336 1330 9432 1346
rect 9336 1194 9366 1330
rect 9564 1296 9594 1594
rect 9792 1426 9822 1594
rect 9872 1532 9902 1594
rect 9872 1502 9930 1532
rect 9726 1410 9822 1426
rect 9726 1376 9742 1410
rect 9776 1376 9822 1410
rect 9726 1360 9822 1376
rect 9498 1280 9594 1296
rect 9498 1246 9514 1280
rect 9548 1246 9594 1280
rect 9498 1230 9594 1246
rect 9564 1194 9594 1230
rect 9792 1194 9822 1360
rect 9900 1344 9930 1502
rect 10128 1426 10158 1594
rect 10208 1532 10238 1594
rect 10208 1502 10266 1532
rect 10062 1410 10158 1426
rect 10062 1376 10078 1410
rect 10112 1376 10158 1410
rect 10062 1360 10158 1376
rect 9900 1328 9996 1344
rect 9900 1294 9946 1328
rect 9980 1294 9996 1328
rect 9900 1278 9996 1294
rect 9900 1194 9930 1278
rect 10128 1194 10158 1360
rect 10236 1344 10266 1502
rect 10504 1426 10534 1594
rect 10438 1410 10534 1426
rect 10438 1376 10454 1410
rect 10488 1376 10534 1410
rect 10438 1360 10534 1376
rect 10236 1328 10332 1344
rect 10236 1294 10282 1328
rect 10316 1294 10332 1328
rect 10236 1278 10332 1294
rect 10236 1194 10266 1278
rect 10504 1194 10534 1360
rect 10772 1296 10802 1594
rect 10852 1532 10882 1594
rect 10852 1502 10910 1532
rect 10706 1280 10802 1296
rect 10706 1246 10722 1280
rect 10756 1246 10802 1280
rect 10706 1230 10802 1246
rect 10772 1194 10802 1230
rect 10880 1396 10910 1502
rect 11108 1396 11138 1594
rect 11188 1532 11218 1594
rect 11188 1502 11246 1532
rect 10880 1380 11138 1396
rect 10880 1346 10990 1380
rect 11024 1346 11138 1380
rect 10880 1330 11138 1346
rect 10880 1194 10910 1330
rect 11108 1194 11138 1330
rect 11216 1396 11246 1502
rect 11216 1380 11312 1396
rect 11216 1346 11262 1380
rect 11296 1346 11312 1380
rect 11216 1330 11312 1346
rect 11216 1194 11246 1330
rect 11444 1296 11474 1594
rect 11672 1426 11702 1594
rect 11752 1532 11782 1594
rect 11752 1502 11810 1532
rect 11606 1410 11702 1426
rect 11606 1376 11622 1410
rect 11656 1376 11702 1410
rect 11606 1360 11702 1376
rect 11378 1280 11474 1296
rect 11378 1246 11394 1280
rect 11428 1246 11474 1280
rect 11378 1230 11474 1246
rect 11444 1194 11474 1230
rect 11672 1194 11702 1360
rect 11780 1344 11810 1502
rect 12008 1426 12038 1594
rect 12088 1532 12118 1594
rect 12088 1502 12146 1532
rect 11942 1410 12038 1426
rect 11942 1376 11958 1410
rect 11992 1376 12038 1410
rect 11942 1360 12038 1376
rect 11780 1328 11876 1344
rect 11780 1294 11826 1328
rect 11860 1294 11876 1328
rect 11780 1278 11876 1294
rect 11780 1194 11810 1278
rect 12008 1194 12038 1360
rect 12116 1344 12146 1502
rect 12116 1328 12212 1344
rect 12116 1294 12162 1328
rect 12196 1294 12212 1328
rect 12344 1296 12374 1594
rect 12424 1532 12454 1594
rect 12424 1502 12482 1532
rect 12116 1278 12212 1294
rect 12278 1280 12374 1296
rect 12116 1194 12146 1278
rect 12278 1246 12294 1280
rect 12328 1246 12374 1280
rect 12278 1230 12374 1246
rect 12344 1194 12374 1230
rect 12452 1396 12482 1502
rect 12680 1396 12710 1594
rect 12760 1532 12790 1594
rect 12760 1502 12818 1532
rect 12452 1380 12710 1396
rect 12452 1346 12562 1380
rect 12596 1346 12710 1380
rect 12452 1330 12710 1346
rect 12452 1194 12482 1330
rect 12680 1194 12710 1330
rect 12788 1396 12818 1502
rect 12788 1380 12884 1396
rect 12788 1346 12834 1380
rect 12868 1346 12884 1380
rect 12788 1330 12884 1346
rect 12788 1194 12818 1330
rect 13016 1296 13046 1594
rect 13244 1426 13274 1594
rect 13324 1532 13354 1594
rect 13324 1502 13382 1532
rect 13178 1410 13274 1426
rect 13178 1376 13194 1410
rect 13228 1376 13274 1410
rect 13178 1360 13274 1376
rect 12950 1280 13046 1296
rect 12950 1246 12966 1280
rect 13000 1246 13046 1280
rect 12950 1230 13046 1246
rect 13016 1194 13046 1230
rect 13244 1194 13274 1360
rect 13352 1344 13382 1502
rect 13580 1426 13610 1594
rect 13660 1532 13690 1594
rect 13660 1502 13718 1532
rect 13514 1410 13610 1426
rect 13514 1376 13530 1410
rect 13564 1376 13610 1410
rect 13514 1360 13610 1376
rect 13352 1328 13448 1344
rect 13352 1294 13398 1328
rect 13432 1294 13448 1328
rect 13352 1278 13448 1294
rect 13352 1194 13382 1278
rect 13580 1194 13610 1360
rect 13688 1344 13718 1502
rect 13688 1328 13784 1344
rect 13688 1294 13734 1328
rect 13768 1294 13784 1328
rect 13688 1278 13784 1294
rect 13688 1194 13718 1278
rect 148 968 178 994
rect 416 968 446 994
rect 524 968 554 994
rect 752 968 782 994
rect 860 968 890 994
rect 1088 968 1118 994
rect 1316 968 1346 994
rect 1424 968 1454 994
rect 1652 968 1682 994
rect 1760 968 1790 994
rect 1988 968 2018 994
rect 2096 968 2126 994
rect 2324 968 2354 994
rect 2432 968 2462 994
rect 2660 968 2690 994
rect 2888 968 2918 994
rect 2996 968 3026 994
rect 3224 968 3254 994
rect 3332 968 3362 994
rect 3600 968 3630 994
rect 3868 968 3898 994
rect 3976 968 4006 994
rect 4204 968 4234 994
rect 4312 968 4342 994
rect 4540 968 4570 994
rect 4768 968 4798 994
rect 4876 968 4906 994
rect 5104 968 5134 994
rect 5212 968 5242 994
rect 5440 968 5470 994
rect 5548 968 5578 994
rect 5776 968 5806 994
rect 5884 968 5914 994
rect 6112 968 6142 994
rect 6340 968 6370 994
rect 6448 968 6478 994
rect 6676 968 6706 994
rect 6784 968 6814 994
rect 7052 968 7082 994
rect 7320 968 7350 994
rect 7428 968 7458 994
rect 7656 968 7686 994
rect 7764 968 7794 994
rect 7992 968 8022 994
rect 8220 968 8250 994
rect 8328 968 8358 994
rect 8556 968 8586 994
rect 8664 968 8694 994
rect 8892 968 8922 994
rect 9000 968 9030 994
rect 9228 968 9258 994
rect 9336 968 9366 994
rect 9564 968 9594 994
rect 9792 968 9822 994
rect 9900 968 9930 994
rect 10128 968 10158 994
rect 10236 968 10266 994
rect 10504 968 10534 994
rect 10772 968 10802 994
rect 10880 968 10910 994
rect 11108 968 11138 994
rect 11216 968 11246 994
rect 11444 968 11474 994
rect 11672 968 11702 994
rect 11780 968 11810 994
rect 12008 968 12038 994
rect 12116 968 12146 994
rect 12344 968 12374 994
rect 12452 968 12482 994
rect 12680 968 12710 994
rect 12788 968 12818 994
rect 13016 968 13046 994
rect 13244 968 13274 994
rect 13352 968 13382 994
rect 13580 968 13610 994
rect 13688 968 13718 994
<< polycont >>
rect 98 1376 132 1410
rect 366 1246 400 1280
rect 634 1346 668 1380
rect 906 1346 940 1380
rect 1266 1376 1300 1410
rect 1038 1246 1072 1280
rect 1602 1376 1636 1410
rect 1470 1294 1504 1328
rect 1806 1294 1840 1328
rect 1938 1246 1972 1280
rect 2206 1346 2240 1380
rect 2478 1346 2512 1380
rect 2838 1376 2872 1410
rect 2610 1246 2644 1280
rect 3174 1376 3208 1410
rect 3042 1294 3076 1328
rect 3550 1376 3584 1410
rect 3378 1294 3412 1328
rect 3818 1246 3852 1280
rect 4086 1346 4120 1380
rect 4358 1346 4392 1380
rect 4718 1376 4752 1410
rect 4490 1246 4524 1280
rect 5054 1376 5088 1410
rect 4922 1294 4956 1328
rect 5258 1294 5292 1328
rect 5390 1246 5424 1280
rect 5658 1346 5692 1380
rect 5930 1346 5964 1380
rect 6290 1376 6324 1410
rect 6062 1246 6096 1280
rect 6626 1376 6660 1410
rect 6494 1294 6528 1328
rect 7002 1376 7036 1410
rect 6830 1294 6864 1328
rect 7270 1246 7304 1280
rect 7538 1346 7572 1380
rect 7810 1346 7844 1380
rect 8170 1376 8204 1410
rect 7942 1246 7976 1280
rect 8506 1376 8540 1410
rect 8374 1294 8408 1328
rect 8710 1294 8744 1328
rect 8842 1246 8876 1280
rect 9110 1346 9144 1380
rect 9382 1346 9416 1380
rect 9742 1376 9776 1410
rect 9514 1246 9548 1280
rect 10078 1376 10112 1410
rect 9946 1294 9980 1328
rect 10454 1376 10488 1410
rect 10282 1294 10316 1328
rect 10722 1246 10756 1280
rect 10990 1346 11024 1380
rect 11262 1346 11296 1380
rect 11622 1376 11656 1410
rect 11394 1246 11428 1280
rect 11958 1376 11992 1410
rect 11826 1294 11860 1328
rect 12162 1294 12196 1328
rect 12294 1246 12328 1280
rect 12562 1346 12596 1380
rect 12834 1346 12868 1380
rect 13194 1376 13228 1410
rect 12966 1246 13000 1280
rect 13530 1376 13564 1410
rect 13398 1294 13432 1328
rect 13734 1294 13768 1328
<< locali >>
rect 4 1804 13862 1824
rect 4 1748 60 1804
rect 266 1748 368 1804
rect 1810 1748 1940 1804
rect 3382 1748 3512 1804
rect 3718 1748 3820 1804
rect 5262 1748 5392 1804
rect 6834 1748 6964 1804
rect 7170 1748 7272 1804
rect 8714 1748 8844 1804
rect 10286 1748 10416 1804
rect 10622 1748 10724 1804
rect 12166 1748 12296 1804
rect 13738 1748 13862 1804
rect 4 1728 13862 1748
rect 76 1678 142 1728
rect 76 1610 92 1678
rect 126 1610 142 1678
rect 76 1594 142 1610
rect 184 1678 250 1694
rect 184 1610 200 1678
rect 234 1610 250 1678
rect 184 1559 250 1610
rect 344 1678 410 1728
rect 344 1610 360 1678
rect 394 1610 410 1678
rect 344 1594 410 1610
rect 532 1678 598 1694
rect 532 1610 548 1678
rect 582 1610 598 1678
rect 184 1493 206 1559
rect 532 1496 598 1610
rect 680 1678 746 1728
rect 680 1610 696 1678
rect 730 1610 746 1678
rect 680 1594 746 1610
rect 868 1678 934 1694
rect 868 1610 884 1678
rect 918 1610 934 1678
rect 868 1580 934 1610
rect 1016 1678 1082 1728
rect 1016 1610 1032 1678
rect 1066 1610 1082 1678
rect 1016 1594 1082 1610
rect 1124 1678 1190 1694
rect 1124 1610 1140 1678
rect 1174 1610 1190 1678
rect 868 1546 884 1580
rect 918 1546 934 1580
rect 868 1496 934 1546
rect 76 1178 142 1194
rect 76 1010 92 1178
rect 126 1010 142 1178
rect 76 960 142 1010
rect 184 1178 250 1493
rect 452 1480 664 1496
rect 452 1446 614 1480
rect 648 1446 664 1480
rect 452 1430 664 1446
rect 788 1430 934 1496
rect 350 1280 416 1296
rect 350 1246 366 1280
rect 400 1246 416 1280
rect 350 1230 416 1246
rect 184 1010 200 1178
rect 234 1010 250 1178
rect 184 994 250 1010
rect 344 1178 410 1194
rect 344 1010 360 1178
rect 394 1010 410 1178
rect 344 960 410 1010
rect 452 1178 518 1430
rect 554 1380 752 1396
rect 554 1346 634 1380
rect 668 1375 752 1380
rect 554 1341 641 1346
rect 675 1341 752 1375
rect 554 1330 752 1341
rect 452 1010 468 1178
rect 502 1010 518 1178
rect 452 994 518 1010
rect 560 1178 626 1194
rect 560 1010 576 1178
rect 610 1010 626 1178
rect 560 960 626 1010
rect 680 1178 746 1194
rect 680 1010 696 1178
rect 730 1010 746 1178
rect 680 960 746 1010
rect 788 1178 854 1430
rect 890 1380 956 1396
rect 890 1346 906 1380
rect 940 1346 956 1380
rect 890 1330 956 1346
rect 1124 1380 1190 1610
rect 1244 1678 1310 1728
rect 1244 1610 1260 1678
rect 1294 1610 1310 1678
rect 1244 1594 1310 1610
rect 1432 1678 1498 1694
rect 1432 1610 1448 1678
rect 1482 1610 1498 1678
rect 1432 1597 1498 1610
rect 1580 1678 1646 1728
rect 1580 1610 1596 1678
rect 1630 1610 1646 1678
rect 1580 1594 1646 1610
rect 1768 1678 1834 1694
rect 1768 1610 1784 1678
rect 1818 1610 1834 1678
rect 1432 1496 1498 1563
rect 1768 1496 1834 1610
rect 1916 1678 1982 1728
rect 1916 1610 1932 1678
rect 1966 1610 1982 1678
rect 1916 1594 1982 1610
rect 2104 1678 2170 1694
rect 2104 1610 2120 1678
rect 2154 1610 2170 1678
rect 2104 1496 2170 1610
rect 2252 1678 2318 1728
rect 2252 1610 2268 1678
rect 2302 1610 2318 1678
rect 2252 1594 2318 1610
rect 2440 1678 2506 1694
rect 2440 1610 2456 1678
rect 2490 1610 2506 1678
rect 2440 1580 2506 1610
rect 2588 1678 2654 1728
rect 2588 1610 2604 1678
rect 2638 1610 2654 1678
rect 2588 1594 2654 1610
rect 2696 1678 2762 1694
rect 2696 1610 2712 1678
rect 2746 1610 2762 1678
rect 2440 1546 2456 1580
rect 2490 1546 2506 1580
rect 2440 1496 2506 1546
rect 1352 1430 1498 1496
rect 1688 1430 1834 1496
rect 2024 1480 2236 1496
rect 2024 1446 2186 1480
rect 2220 1446 2236 1480
rect 2024 1430 2236 1446
rect 2360 1430 2506 1496
rect 1124 1346 1140 1380
rect 1174 1346 1190 1380
rect 1250 1410 1316 1426
rect 1250 1376 1266 1410
rect 1300 1376 1316 1410
rect 1250 1360 1316 1376
rect 1352 1410 1418 1430
rect 1352 1376 1368 1410
rect 1402 1376 1418 1410
rect 1022 1280 1088 1296
rect 1022 1246 1038 1280
rect 1072 1246 1088 1280
rect 1022 1230 1088 1246
rect 788 1010 804 1178
rect 838 1010 854 1178
rect 788 994 854 1010
rect 896 1178 962 1194
rect 896 1010 912 1178
rect 946 1010 962 1178
rect 896 960 962 1010
rect 1016 1178 1082 1194
rect 1016 1010 1032 1178
rect 1066 1010 1082 1178
rect 1016 960 1082 1010
rect 1124 1178 1190 1346
rect 1124 1010 1140 1178
rect 1174 1010 1190 1178
rect 1124 994 1190 1010
rect 1244 1178 1310 1194
rect 1244 1010 1260 1178
rect 1294 1010 1310 1178
rect 1244 960 1310 1010
rect 1352 1178 1418 1376
rect 1586 1410 1652 1426
rect 1586 1376 1602 1410
rect 1636 1376 1652 1410
rect 1586 1360 1652 1376
rect 1454 1328 1520 1344
rect 1454 1294 1470 1328
rect 1504 1294 1520 1328
rect 1454 1278 1520 1294
rect 1688 1328 1754 1430
rect 1688 1294 1704 1328
rect 1738 1294 1754 1328
rect 1352 1010 1368 1178
rect 1402 1010 1418 1178
rect 1352 994 1418 1010
rect 1460 1178 1526 1194
rect 1460 1010 1476 1178
rect 1510 1010 1526 1178
rect 1460 960 1526 1010
rect 1580 1178 1646 1194
rect 1580 1010 1596 1178
rect 1630 1010 1646 1178
rect 1580 960 1646 1010
rect 1688 1178 1754 1294
rect 1790 1328 1856 1344
rect 1790 1294 1806 1328
rect 1840 1294 1856 1328
rect 1790 1278 1856 1294
rect 1922 1280 1988 1296
rect 1922 1246 1938 1280
rect 1972 1246 1988 1280
rect 1922 1230 1988 1246
rect 1688 1010 1704 1178
rect 1738 1010 1754 1178
rect 1688 994 1754 1010
rect 1796 1178 1862 1194
rect 1796 1010 1812 1178
rect 1846 1010 1862 1178
rect 1796 960 1862 1010
rect 1916 1178 1982 1194
rect 1916 1010 1932 1178
rect 1966 1010 1982 1178
rect 1916 960 1982 1010
rect 2024 1178 2090 1430
rect 2126 1381 2324 1396
rect 2126 1380 2209 1381
rect 2126 1346 2206 1380
rect 2243 1347 2324 1381
rect 2240 1346 2324 1347
rect 2126 1330 2324 1346
rect 2024 1010 2040 1178
rect 2074 1010 2090 1178
rect 2024 994 2090 1010
rect 2132 1178 2198 1194
rect 2132 1010 2148 1178
rect 2182 1010 2198 1178
rect 2132 960 2198 1010
rect 2252 1178 2318 1194
rect 2252 1010 2268 1178
rect 2302 1010 2318 1178
rect 2252 960 2318 1010
rect 2360 1178 2426 1430
rect 2462 1380 2528 1396
rect 2462 1346 2478 1380
rect 2512 1346 2528 1380
rect 2462 1330 2528 1346
rect 2696 1380 2762 1610
rect 2816 1678 2882 1728
rect 2816 1610 2832 1678
rect 2866 1610 2882 1678
rect 2816 1594 2882 1610
rect 3004 1678 3070 1694
rect 3004 1610 3020 1678
rect 3054 1610 3070 1678
rect 3004 1496 3070 1610
rect 3152 1678 3218 1728
rect 3152 1610 3168 1678
rect 3202 1610 3218 1678
rect 3152 1594 3218 1610
rect 3340 1678 3406 1694
rect 3340 1610 3356 1678
rect 3390 1610 3406 1678
rect 3340 1496 3406 1610
rect 3528 1678 3594 1728
rect 3528 1610 3544 1678
rect 3578 1610 3594 1678
rect 3528 1594 3594 1610
rect 3636 1678 3702 1694
rect 3636 1610 3652 1678
rect 3686 1610 3702 1678
rect 2924 1430 3070 1496
rect 3260 1430 3406 1496
rect 3636 1559 3702 1610
rect 3796 1678 3862 1728
rect 3796 1610 3812 1678
rect 3846 1610 3862 1678
rect 3796 1594 3862 1610
rect 3984 1678 4050 1694
rect 3984 1610 4000 1678
rect 4034 1610 4050 1678
rect 3636 1493 3658 1559
rect 3984 1496 4050 1610
rect 4132 1678 4198 1728
rect 4132 1610 4148 1678
rect 4182 1610 4198 1678
rect 4132 1594 4198 1610
rect 4320 1678 4386 1694
rect 4320 1610 4336 1678
rect 4370 1610 4386 1678
rect 4320 1580 4386 1610
rect 4468 1678 4534 1728
rect 4468 1610 4484 1678
rect 4518 1610 4534 1678
rect 4468 1594 4534 1610
rect 4576 1678 4642 1694
rect 4576 1610 4592 1678
rect 4626 1610 4642 1678
rect 4320 1546 4336 1580
rect 4370 1546 4386 1580
rect 4320 1496 4386 1546
rect 2696 1346 2712 1380
rect 2746 1346 2762 1380
rect 2822 1410 2888 1426
rect 2822 1376 2838 1410
rect 2872 1376 2888 1410
rect 2822 1360 2888 1376
rect 2924 1410 2990 1430
rect 2924 1376 2940 1410
rect 2974 1376 2990 1410
rect 2594 1280 2660 1296
rect 2594 1246 2610 1280
rect 2644 1246 2660 1280
rect 2594 1230 2660 1246
rect 2360 1010 2376 1178
rect 2410 1010 2426 1178
rect 2360 994 2426 1010
rect 2468 1178 2534 1194
rect 2468 1010 2484 1178
rect 2518 1010 2534 1178
rect 2468 960 2534 1010
rect 2588 1178 2654 1194
rect 2588 1010 2604 1178
rect 2638 1010 2654 1178
rect 2588 960 2654 1010
rect 2696 1178 2762 1346
rect 2696 1010 2712 1178
rect 2746 1010 2762 1178
rect 2696 994 2762 1010
rect 2816 1178 2882 1194
rect 2816 1010 2832 1178
rect 2866 1010 2882 1178
rect 2816 960 2882 1010
rect 2924 1178 2990 1376
rect 3158 1410 3224 1426
rect 3158 1376 3174 1410
rect 3208 1376 3224 1410
rect 3158 1360 3224 1376
rect 3026 1328 3092 1344
rect 3026 1294 3042 1328
rect 3076 1294 3092 1328
rect 3026 1278 3092 1294
rect 3260 1328 3326 1430
rect 3260 1294 3276 1328
rect 3310 1294 3326 1328
rect 2924 1010 2940 1178
rect 2974 1010 2990 1178
rect 2924 994 2990 1010
rect 3032 1178 3098 1194
rect 3032 1010 3048 1178
rect 3082 1010 3098 1178
rect 3032 960 3098 1010
rect 3152 1178 3218 1194
rect 3152 1010 3168 1178
rect 3202 1010 3218 1178
rect 3152 960 3218 1010
rect 3260 1178 3326 1294
rect 3362 1328 3428 1344
rect 3362 1294 3378 1328
rect 3412 1294 3428 1328
rect 3362 1278 3428 1294
rect 3260 1010 3276 1178
rect 3310 1010 3326 1178
rect 3260 994 3326 1010
rect 3368 1178 3434 1194
rect 3368 1010 3384 1178
rect 3418 1010 3434 1178
rect 3368 960 3434 1010
rect 3528 1178 3594 1194
rect 3528 1010 3544 1178
rect 3578 1010 3594 1178
rect 3528 960 3594 1010
rect 3636 1178 3702 1493
rect 3904 1480 4116 1496
rect 3904 1446 4066 1480
rect 4100 1446 4116 1480
rect 3904 1430 4116 1446
rect 4240 1430 4386 1496
rect 3802 1280 3868 1296
rect 3802 1246 3818 1280
rect 3852 1246 3868 1280
rect 3802 1230 3868 1246
rect 3636 1010 3652 1178
rect 3686 1010 3702 1178
rect 3636 994 3702 1010
rect 3796 1178 3862 1194
rect 3796 1010 3812 1178
rect 3846 1010 3862 1178
rect 3796 960 3862 1010
rect 3904 1178 3970 1430
rect 4006 1380 4204 1396
rect 4006 1346 4086 1380
rect 4120 1375 4204 1380
rect 4006 1341 4093 1346
rect 4127 1341 4204 1375
rect 4006 1330 4204 1341
rect 3904 1010 3920 1178
rect 3954 1010 3970 1178
rect 3904 994 3970 1010
rect 4012 1178 4078 1194
rect 4012 1010 4028 1178
rect 4062 1010 4078 1178
rect 4012 960 4078 1010
rect 4132 1178 4198 1194
rect 4132 1010 4148 1178
rect 4182 1010 4198 1178
rect 4132 960 4198 1010
rect 4240 1178 4306 1430
rect 4342 1380 4408 1396
rect 4342 1346 4358 1380
rect 4392 1346 4408 1380
rect 4342 1330 4408 1346
rect 4576 1380 4642 1610
rect 4696 1678 4762 1728
rect 4696 1610 4712 1678
rect 4746 1610 4762 1678
rect 4696 1594 4762 1610
rect 4884 1678 4950 1694
rect 4884 1610 4900 1678
rect 4934 1610 4950 1678
rect 4884 1597 4950 1610
rect 5032 1678 5098 1728
rect 5032 1610 5048 1678
rect 5082 1610 5098 1678
rect 5032 1594 5098 1610
rect 5220 1678 5286 1694
rect 5220 1610 5236 1678
rect 5270 1610 5286 1678
rect 4884 1496 4950 1563
rect 5220 1496 5286 1610
rect 5368 1678 5434 1728
rect 5368 1610 5384 1678
rect 5418 1610 5434 1678
rect 5368 1594 5434 1610
rect 5556 1678 5622 1694
rect 5556 1610 5572 1678
rect 5606 1610 5622 1678
rect 5556 1496 5622 1610
rect 5704 1678 5770 1728
rect 5704 1610 5720 1678
rect 5754 1610 5770 1678
rect 5704 1594 5770 1610
rect 5892 1678 5958 1694
rect 5892 1610 5908 1678
rect 5942 1610 5958 1678
rect 5892 1580 5958 1610
rect 6040 1678 6106 1728
rect 6040 1610 6056 1678
rect 6090 1610 6106 1678
rect 6040 1594 6106 1610
rect 6148 1678 6214 1694
rect 6148 1610 6164 1678
rect 6198 1610 6214 1678
rect 5892 1546 5908 1580
rect 5942 1546 5958 1580
rect 5892 1496 5958 1546
rect 4804 1430 4950 1496
rect 5140 1430 5286 1496
rect 5476 1480 5688 1496
rect 5476 1446 5638 1480
rect 5672 1446 5688 1480
rect 5476 1430 5688 1446
rect 5812 1430 5958 1496
rect 4576 1346 4592 1380
rect 4626 1346 4642 1380
rect 4702 1410 4768 1426
rect 4702 1376 4718 1410
rect 4752 1376 4768 1410
rect 4702 1360 4768 1376
rect 4804 1410 4870 1430
rect 4804 1376 4820 1410
rect 4854 1376 4870 1410
rect 4474 1280 4540 1296
rect 4474 1246 4490 1280
rect 4524 1246 4540 1280
rect 4474 1230 4540 1246
rect 4240 1010 4256 1178
rect 4290 1010 4306 1178
rect 4240 994 4306 1010
rect 4348 1178 4414 1194
rect 4348 1010 4364 1178
rect 4398 1010 4414 1178
rect 4348 960 4414 1010
rect 4468 1178 4534 1194
rect 4468 1010 4484 1178
rect 4518 1010 4534 1178
rect 4468 960 4534 1010
rect 4576 1178 4642 1346
rect 4576 1010 4592 1178
rect 4626 1010 4642 1178
rect 4576 994 4642 1010
rect 4696 1178 4762 1194
rect 4696 1010 4712 1178
rect 4746 1010 4762 1178
rect 4696 960 4762 1010
rect 4804 1178 4870 1376
rect 5038 1410 5104 1426
rect 5038 1376 5054 1410
rect 5088 1376 5104 1410
rect 5038 1360 5104 1376
rect 4906 1328 4972 1344
rect 4906 1294 4922 1328
rect 4956 1294 4972 1328
rect 4906 1278 4972 1294
rect 5140 1328 5206 1430
rect 5140 1294 5156 1328
rect 5190 1294 5206 1328
rect 4804 1010 4820 1178
rect 4854 1010 4870 1178
rect 4804 994 4870 1010
rect 4912 1178 4978 1194
rect 4912 1010 4928 1178
rect 4962 1010 4978 1178
rect 4912 960 4978 1010
rect 5032 1178 5098 1194
rect 5032 1010 5048 1178
rect 5082 1010 5098 1178
rect 5032 960 5098 1010
rect 5140 1178 5206 1294
rect 5242 1328 5308 1344
rect 5242 1294 5258 1328
rect 5292 1294 5308 1328
rect 5242 1278 5308 1294
rect 5374 1280 5440 1296
rect 5374 1246 5390 1280
rect 5424 1246 5440 1280
rect 5374 1230 5440 1246
rect 5140 1010 5156 1178
rect 5190 1010 5206 1178
rect 5140 994 5206 1010
rect 5248 1178 5314 1194
rect 5248 1010 5264 1178
rect 5298 1010 5314 1178
rect 5248 960 5314 1010
rect 5368 1178 5434 1194
rect 5368 1010 5384 1178
rect 5418 1010 5434 1178
rect 5368 960 5434 1010
rect 5476 1178 5542 1430
rect 5578 1381 5776 1396
rect 5578 1380 5661 1381
rect 5578 1346 5658 1380
rect 5695 1347 5776 1381
rect 5692 1346 5776 1347
rect 5578 1330 5776 1346
rect 5476 1010 5492 1178
rect 5526 1010 5542 1178
rect 5476 994 5542 1010
rect 5584 1178 5650 1194
rect 5584 1010 5600 1178
rect 5634 1010 5650 1178
rect 5584 960 5650 1010
rect 5704 1178 5770 1194
rect 5704 1010 5720 1178
rect 5754 1010 5770 1178
rect 5704 960 5770 1010
rect 5812 1178 5878 1430
rect 5914 1380 5980 1396
rect 5914 1346 5930 1380
rect 5964 1346 5980 1380
rect 5914 1330 5980 1346
rect 6148 1380 6214 1610
rect 6268 1678 6334 1728
rect 6268 1610 6284 1678
rect 6318 1610 6334 1678
rect 6268 1594 6334 1610
rect 6456 1678 6522 1694
rect 6456 1610 6472 1678
rect 6506 1610 6522 1678
rect 6456 1496 6522 1610
rect 6604 1678 6670 1728
rect 6604 1610 6620 1678
rect 6654 1610 6670 1678
rect 6604 1594 6670 1610
rect 6792 1678 6858 1694
rect 6792 1610 6808 1678
rect 6842 1610 6858 1678
rect 6792 1496 6858 1610
rect 6980 1678 7046 1728
rect 6980 1610 6996 1678
rect 7030 1610 7046 1678
rect 6980 1594 7046 1610
rect 7088 1678 7154 1694
rect 7088 1610 7104 1678
rect 7138 1610 7154 1678
rect 6376 1430 6522 1496
rect 6712 1430 6858 1496
rect 7088 1559 7154 1610
rect 7248 1678 7314 1728
rect 7248 1610 7264 1678
rect 7298 1610 7314 1678
rect 7248 1594 7314 1610
rect 7436 1678 7502 1694
rect 7436 1610 7452 1678
rect 7486 1610 7502 1678
rect 7088 1493 7110 1559
rect 7436 1496 7502 1610
rect 7584 1678 7650 1728
rect 7584 1610 7600 1678
rect 7634 1610 7650 1678
rect 7584 1594 7650 1610
rect 7772 1678 7838 1694
rect 7772 1610 7788 1678
rect 7822 1610 7838 1678
rect 7772 1580 7838 1610
rect 7920 1678 7986 1728
rect 7920 1610 7936 1678
rect 7970 1610 7986 1678
rect 7920 1594 7986 1610
rect 8028 1678 8094 1694
rect 8028 1610 8044 1678
rect 8078 1610 8094 1678
rect 7772 1546 7788 1580
rect 7822 1546 7838 1580
rect 7772 1496 7838 1546
rect 6148 1346 6164 1380
rect 6198 1346 6214 1380
rect 6274 1410 6340 1426
rect 6274 1376 6290 1410
rect 6324 1376 6340 1410
rect 6274 1360 6340 1376
rect 6376 1410 6442 1430
rect 6376 1376 6392 1410
rect 6426 1376 6442 1410
rect 6046 1280 6112 1296
rect 6046 1246 6062 1280
rect 6096 1246 6112 1280
rect 6046 1230 6112 1246
rect 5812 1010 5828 1178
rect 5862 1010 5878 1178
rect 5812 994 5878 1010
rect 5920 1178 5986 1194
rect 5920 1010 5936 1178
rect 5970 1010 5986 1178
rect 5920 960 5986 1010
rect 6040 1178 6106 1194
rect 6040 1010 6056 1178
rect 6090 1010 6106 1178
rect 6040 960 6106 1010
rect 6148 1178 6214 1346
rect 6148 1010 6164 1178
rect 6198 1010 6214 1178
rect 6148 994 6214 1010
rect 6268 1178 6334 1194
rect 6268 1010 6284 1178
rect 6318 1010 6334 1178
rect 6268 960 6334 1010
rect 6376 1178 6442 1376
rect 6610 1410 6676 1426
rect 6610 1376 6626 1410
rect 6660 1376 6676 1410
rect 6610 1360 6676 1376
rect 6478 1328 6544 1344
rect 6478 1294 6494 1328
rect 6528 1294 6544 1328
rect 6478 1278 6544 1294
rect 6712 1328 6778 1430
rect 6712 1294 6728 1328
rect 6762 1294 6778 1328
rect 6376 1010 6392 1178
rect 6426 1010 6442 1178
rect 6376 994 6442 1010
rect 6484 1178 6550 1194
rect 6484 1010 6500 1178
rect 6534 1010 6550 1178
rect 6484 960 6550 1010
rect 6604 1178 6670 1194
rect 6604 1010 6620 1178
rect 6654 1010 6670 1178
rect 6604 960 6670 1010
rect 6712 1178 6778 1294
rect 6814 1328 6880 1344
rect 6814 1294 6830 1328
rect 6864 1294 6880 1328
rect 6814 1278 6880 1294
rect 6712 1010 6728 1178
rect 6762 1010 6778 1178
rect 6712 994 6778 1010
rect 6820 1178 6886 1194
rect 6820 1010 6836 1178
rect 6870 1010 6886 1178
rect 6820 960 6886 1010
rect 6980 1178 7046 1194
rect 6980 1010 6996 1178
rect 7030 1010 7046 1178
rect 6980 960 7046 1010
rect 7088 1178 7154 1493
rect 7356 1480 7568 1496
rect 7356 1446 7518 1480
rect 7552 1446 7568 1480
rect 7356 1430 7568 1446
rect 7692 1430 7838 1496
rect 7254 1280 7320 1296
rect 7254 1246 7270 1280
rect 7304 1246 7320 1280
rect 7254 1230 7320 1246
rect 7088 1010 7104 1178
rect 7138 1010 7154 1178
rect 7088 994 7154 1010
rect 7248 1178 7314 1194
rect 7248 1010 7264 1178
rect 7298 1010 7314 1178
rect 7248 960 7314 1010
rect 7356 1178 7422 1430
rect 7458 1380 7656 1396
rect 7458 1346 7538 1380
rect 7572 1375 7656 1380
rect 7458 1341 7545 1346
rect 7579 1341 7656 1375
rect 7458 1330 7656 1341
rect 7356 1010 7372 1178
rect 7406 1010 7422 1178
rect 7356 994 7422 1010
rect 7464 1178 7530 1194
rect 7464 1010 7480 1178
rect 7514 1010 7530 1178
rect 7464 960 7530 1010
rect 7584 1178 7650 1194
rect 7584 1010 7600 1178
rect 7634 1010 7650 1178
rect 7584 960 7650 1010
rect 7692 1178 7758 1430
rect 7794 1380 7860 1396
rect 7794 1346 7810 1380
rect 7844 1346 7860 1380
rect 7794 1330 7860 1346
rect 8028 1380 8094 1610
rect 8148 1678 8214 1728
rect 8148 1610 8164 1678
rect 8198 1610 8214 1678
rect 8148 1594 8214 1610
rect 8336 1678 8402 1694
rect 8336 1610 8352 1678
rect 8386 1610 8402 1678
rect 8336 1597 8402 1610
rect 8484 1678 8550 1728
rect 8484 1610 8500 1678
rect 8534 1610 8550 1678
rect 8484 1594 8550 1610
rect 8672 1678 8738 1694
rect 8672 1610 8688 1678
rect 8722 1610 8738 1678
rect 8336 1496 8402 1563
rect 8672 1496 8738 1610
rect 8820 1678 8886 1728
rect 8820 1610 8836 1678
rect 8870 1610 8886 1678
rect 8820 1594 8886 1610
rect 9008 1678 9074 1694
rect 9008 1610 9024 1678
rect 9058 1610 9074 1678
rect 9008 1496 9074 1610
rect 9156 1678 9222 1728
rect 9156 1610 9172 1678
rect 9206 1610 9222 1678
rect 9156 1594 9222 1610
rect 9344 1678 9410 1694
rect 9344 1610 9360 1678
rect 9394 1610 9410 1678
rect 9344 1580 9410 1610
rect 9492 1678 9558 1728
rect 9492 1610 9508 1678
rect 9542 1610 9558 1678
rect 9492 1594 9558 1610
rect 9600 1678 9666 1694
rect 9600 1610 9616 1678
rect 9650 1610 9666 1678
rect 9344 1546 9360 1580
rect 9394 1546 9410 1580
rect 9344 1496 9410 1546
rect 8256 1430 8402 1496
rect 8592 1430 8738 1496
rect 8928 1480 9140 1496
rect 8928 1446 9090 1480
rect 9124 1446 9140 1480
rect 8928 1430 9140 1446
rect 9264 1430 9410 1496
rect 8028 1346 8044 1380
rect 8078 1346 8094 1380
rect 8154 1410 8220 1426
rect 8154 1376 8170 1410
rect 8204 1376 8220 1410
rect 8154 1360 8220 1376
rect 8256 1410 8322 1430
rect 8256 1376 8272 1410
rect 8306 1376 8322 1410
rect 7926 1280 7992 1296
rect 7926 1246 7942 1280
rect 7976 1246 7992 1280
rect 7926 1230 7992 1246
rect 7692 1010 7708 1178
rect 7742 1010 7758 1178
rect 7692 994 7758 1010
rect 7800 1178 7866 1194
rect 7800 1010 7816 1178
rect 7850 1010 7866 1178
rect 7800 960 7866 1010
rect 7920 1178 7986 1194
rect 7920 1010 7936 1178
rect 7970 1010 7986 1178
rect 7920 960 7986 1010
rect 8028 1178 8094 1346
rect 8028 1010 8044 1178
rect 8078 1010 8094 1178
rect 8028 994 8094 1010
rect 8148 1178 8214 1194
rect 8148 1010 8164 1178
rect 8198 1010 8214 1178
rect 8148 960 8214 1010
rect 8256 1178 8322 1376
rect 8490 1410 8556 1426
rect 8490 1376 8506 1410
rect 8540 1376 8556 1410
rect 8490 1360 8556 1376
rect 8358 1328 8424 1344
rect 8358 1294 8374 1328
rect 8408 1294 8424 1328
rect 8358 1278 8424 1294
rect 8592 1328 8658 1430
rect 8592 1294 8608 1328
rect 8642 1294 8658 1328
rect 8256 1010 8272 1178
rect 8306 1010 8322 1178
rect 8256 994 8322 1010
rect 8364 1178 8430 1194
rect 8364 1010 8380 1178
rect 8414 1010 8430 1178
rect 8364 960 8430 1010
rect 8484 1178 8550 1194
rect 8484 1010 8500 1178
rect 8534 1010 8550 1178
rect 8484 960 8550 1010
rect 8592 1178 8658 1294
rect 8694 1328 8760 1344
rect 8694 1294 8710 1328
rect 8744 1294 8760 1328
rect 8694 1278 8760 1294
rect 8826 1280 8892 1296
rect 8826 1246 8842 1280
rect 8876 1246 8892 1280
rect 8826 1230 8892 1246
rect 8592 1010 8608 1178
rect 8642 1010 8658 1178
rect 8592 994 8658 1010
rect 8700 1178 8766 1194
rect 8700 1010 8716 1178
rect 8750 1010 8766 1178
rect 8700 960 8766 1010
rect 8820 1178 8886 1194
rect 8820 1010 8836 1178
rect 8870 1010 8886 1178
rect 8820 960 8886 1010
rect 8928 1178 8994 1430
rect 9030 1381 9228 1396
rect 9030 1380 9113 1381
rect 9030 1346 9110 1380
rect 9147 1347 9228 1381
rect 9144 1346 9228 1347
rect 9030 1330 9228 1346
rect 8928 1010 8944 1178
rect 8978 1010 8994 1178
rect 8928 994 8994 1010
rect 9036 1178 9102 1194
rect 9036 1010 9052 1178
rect 9086 1010 9102 1178
rect 9036 960 9102 1010
rect 9156 1178 9222 1194
rect 9156 1010 9172 1178
rect 9206 1010 9222 1178
rect 9156 960 9222 1010
rect 9264 1178 9330 1430
rect 9366 1380 9432 1396
rect 9366 1346 9382 1380
rect 9416 1346 9432 1380
rect 9366 1330 9432 1346
rect 9600 1380 9666 1610
rect 9720 1678 9786 1728
rect 9720 1610 9736 1678
rect 9770 1610 9786 1678
rect 9720 1594 9786 1610
rect 9908 1678 9974 1694
rect 9908 1610 9924 1678
rect 9958 1610 9974 1678
rect 9908 1496 9974 1610
rect 10056 1678 10122 1728
rect 10056 1610 10072 1678
rect 10106 1610 10122 1678
rect 10056 1594 10122 1610
rect 10244 1678 10310 1694
rect 10244 1610 10260 1678
rect 10294 1610 10310 1678
rect 10244 1496 10310 1610
rect 10432 1678 10498 1728
rect 10432 1610 10448 1678
rect 10482 1610 10498 1678
rect 10432 1594 10498 1610
rect 10540 1678 10606 1694
rect 10540 1610 10556 1678
rect 10590 1610 10606 1678
rect 9828 1430 9974 1496
rect 10164 1430 10310 1496
rect 10540 1559 10606 1610
rect 10700 1678 10766 1728
rect 10700 1610 10716 1678
rect 10750 1610 10766 1678
rect 10700 1594 10766 1610
rect 10888 1678 10954 1694
rect 10888 1610 10904 1678
rect 10938 1610 10954 1678
rect 10540 1493 10562 1559
rect 10888 1496 10954 1610
rect 11036 1678 11102 1728
rect 11036 1610 11052 1678
rect 11086 1610 11102 1678
rect 11036 1594 11102 1610
rect 11224 1678 11290 1694
rect 11224 1610 11240 1678
rect 11274 1610 11290 1678
rect 11224 1580 11290 1610
rect 11372 1678 11438 1728
rect 11372 1610 11388 1678
rect 11422 1610 11438 1678
rect 11372 1594 11438 1610
rect 11480 1678 11546 1694
rect 11480 1610 11496 1678
rect 11530 1610 11546 1678
rect 11224 1546 11240 1580
rect 11274 1546 11290 1580
rect 11224 1496 11290 1546
rect 9600 1346 9616 1380
rect 9650 1346 9666 1380
rect 9726 1410 9792 1426
rect 9726 1376 9742 1410
rect 9776 1376 9792 1410
rect 9726 1360 9792 1376
rect 9828 1410 9894 1430
rect 9828 1376 9844 1410
rect 9878 1376 9894 1410
rect 9498 1280 9564 1296
rect 9498 1246 9514 1280
rect 9548 1246 9564 1280
rect 9498 1230 9564 1246
rect 9264 1010 9280 1178
rect 9314 1010 9330 1178
rect 9264 994 9330 1010
rect 9372 1178 9438 1194
rect 9372 1010 9388 1178
rect 9422 1010 9438 1178
rect 9372 960 9438 1010
rect 9492 1178 9558 1194
rect 9492 1010 9508 1178
rect 9542 1010 9558 1178
rect 9492 960 9558 1010
rect 9600 1178 9666 1346
rect 9600 1010 9616 1178
rect 9650 1010 9666 1178
rect 9600 994 9666 1010
rect 9720 1178 9786 1194
rect 9720 1010 9736 1178
rect 9770 1010 9786 1178
rect 9720 960 9786 1010
rect 9828 1178 9894 1376
rect 10062 1410 10128 1426
rect 10062 1376 10078 1410
rect 10112 1376 10128 1410
rect 10062 1360 10128 1376
rect 9930 1328 9996 1344
rect 9930 1294 9946 1328
rect 9980 1294 9996 1328
rect 9930 1278 9996 1294
rect 10164 1328 10230 1430
rect 10164 1294 10180 1328
rect 10214 1294 10230 1328
rect 9828 1010 9844 1178
rect 9878 1010 9894 1178
rect 9828 994 9894 1010
rect 9936 1178 10002 1194
rect 9936 1010 9952 1178
rect 9986 1010 10002 1178
rect 9936 960 10002 1010
rect 10056 1178 10122 1194
rect 10056 1010 10072 1178
rect 10106 1010 10122 1178
rect 10056 960 10122 1010
rect 10164 1178 10230 1294
rect 10266 1328 10332 1344
rect 10266 1294 10282 1328
rect 10316 1294 10332 1328
rect 10266 1278 10332 1294
rect 10164 1010 10180 1178
rect 10214 1010 10230 1178
rect 10164 994 10230 1010
rect 10272 1178 10338 1194
rect 10272 1010 10288 1178
rect 10322 1010 10338 1178
rect 10272 960 10338 1010
rect 10432 1178 10498 1194
rect 10432 1010 10448 1178
rect 10482 1010 10498 1178
rect 10432 960 10498 1010
rect 10540 1178 10606 1493
rect 10808 1480 11020 1496
rect 10808 1446 10970 1480
rect 11004 1446 11020 1480
rect 10808 1430 11020 1446
rect 11144 1430 11290 1496
rect 10706 1280 10772 1296
rect 10706 1246 10722 1280
rect 10756 1246 10772 1280
rect 10706 1230 10772 1246
rect 10540 1010 10556 1178
rect 10590 1010 10606 1178
rect 10540 994 10606 1010
rect 10700 1178 10766 1194
rect 10700 1010 10716 1178
rect 10750 1010 10766 1178
rect 10700 960 10766 1010
rect 10808 1178 10874 1430
rect 10910 1380 11108 1396
rect 10910 1346 10990 1380
rect 11024 1375 11108 1380
rect 10910 1341 10997 1346
rect 11031 1341 11108 1375
rect 10910 1330 11108 1341
rect 10808 1010 10824 1178
rect 10858 1010 10874 1178
rect 10808 994 10874 1010
rect 10916 1178 10982 1194
rect 10916 1010 10932 1178
rect 10966 1010 10982 1178
rect 10916 960 10982 1010
rect 11036 1178 11102 1194
rect 11036 1010 11052 1178
rect 11086 1010 11102 1178
rect 11036 960 11102 1010
rect 11144 1178 11210 1430
rect 11246 1380 11312 1396
rect 11246 1346 11262 1380
rect 11296 1346 11312 1380
rect 11246 1330 11312 1346
rect 11480 1380 11546 1610
rect 11600 1678 11666 1728
rect 11600 1610 11616 1678
rect 11650 1610 11666 1678
rect 11600 1594 11666 1610
rect 11788 1678 11854 1694
rect 11788 1610 11804 1678
rect 11838 1610 11854 1678
rect 11788 1597 11854 1610
rect 11936 1678 12002 1728
rect 11936 1610 11952 1678
rect 11986 1610 12002 1678
rect 11936 1594 12002 1610
rect 12124 1678 12190 1694
rect 12124 1610 12140 1678
rect 12174 1610 12190 1678
rect 11788 1496 11854 1563
rect 12124 1496 12190 1610
rect 12272 1678 12338 1728
rect 12272 1610 12288 1678
rect 12322 1610 12338 1678
rect 12272 1594 12338 1610
rect 12460 1678 12526 1694
rect 12460 1610 12476 1678
rect 12510 1610 12526 1678
rect 12460 1496 12526 1610
rect 12608 1678 12674 1728
rect 12608 1610 12624 1678
rect 12658 1610 12674 1678
rect 12608 1594 12674 1610
rect 12796 1678 12862 1694
rect 12796 1610 12812 1678
rect 12846 1610 12862 1678
rect 12796 1580 12862 1610
rect 12944 1678 13010 1728
rect 12944 1610 12960 1678
rect 12994 1610 13010 1678
rect 12944 1594 13010 1610
rect 13052 1678 13118 1694
rect 13052 1610 13068 1678
rect 13102 1610 13118 1678
rect 12796 1546 12812 1580
rect 12846 1546 12862 1580
rect 12796 1496 12862 1546
rect 11708 1430 11854 1496
rect 12044 1430 12190 1496
rect 12380 1480 12592 1496
rect 12380 1446 12542 1480
rect 12576 1446 12592 1480
rect 12380 1430 12592 1446
rect 12716 1430 12862 1496
rect 11480 1346 11496 1380
rect 11530 1346 11546 1380
rect 11606 1410 11672 1426
rect 11606 1376 11622 1410
rect 11656 1376 11672 1410
rect 11606 1360 11672 1376
rect 11708 1410 11774 1430
rect 11708 1376 11724 1410
rect 11758 1376 11774 1410
rect 11378 1280 11444 1296
rect 11378 1246 11394 1280
rect 11428 1246 11444 1280
rect 11378 1230 11444 1246
rect 11144 1010 11160 1178
rect 11194 1010 11210 1178
rect 11144 994 11210 1010
rect 11252 1178 11318 1194
rect 11252 1010 11268 1178
rect 11302 1010 11318 1178
rect 11252 960 11318 1010
rect 11372 1178 11438 1194
rect 11372 1010 11388 1178
rect 11422 1010 11438 1178
rect 11372 960 11438 1010
rect 11480 1178 11546 1346
rect 11480 1010 11496 1178
rect 11530 1010 11546 1178
rect 11480 994 11546 1010
rect 11600 1178 11666 1194
rect 11600 1010 11616 1178
rect 11650 1010 11666 1178
rect 11600 960 11666 1010
rect 11708 1178 11774 1376
rect 11942 1410 12008 1426
rect 11942 1376 11958 1410
rect 11992 1376 12008 1410
rect 11942 1360 12008 1376
rect 11810 1328 11876 1344
rect 11810 1294 11826 1328
rect 11860 1294 11876 1328
rect 11810 1278 11876 1294
rect 12044 1328 12110 1430
rect 12044 1294 12060 1328
rect 12094 1294 12110 1328
rect 11708 1010 11724 1178
rect 11758 1010 11774 1178
rect 11708 994 11774 1010
rect 11816 1178 11882 1194
rect 11816 1010 11832 1178
rect 11866 1010 11882 1178
rect 11816 960 11882 1010
rect 11936 1178 12002 1194
rect 11936 1010 11952 1178
rect 11986 1010 12002 1178
rect 11936 960 12002 1010
rect 12044 1178 12110 1294
rect 12146 1328 12212 1344
rect 12146 1294 12162 1328
rect 12196 1294 12212 1328
rect 12146 1278 12212 1294
rect 12278 1280 12344 1296
rect 12278 1246 12294 1280
rect 12328 1246 12344 1280
rect 12278 1230 12344 1246
rect 12044 1010 12060 1178
rect 12094 1010 12110 1178
rect 12044 994 12110 1010
rect 12152 1178 12218 1194
rect 12152 1010 12168 1178
rect 12202 1010 12218 1178
rect 12152 960 12218 1010
rect 12272 1178 12338 1194
rect 12272 1010 12288 1178
rect 12322 1010 12338 1178
rect 12272 960 12338 1010
rect 12380 1178 12446 1430
rect 12482 1381 12680 1396
rect 12482 1380 12565 1381
rect 12482 1346 12562 1380
rect 12599 1347 12680 1381
rect 12596 1346 12680 1347
rect 12482 1330 12680 1346
rect 12380 1010 12396 1178
rect 12430 1010 12446 1178
rect 12380 994 12446 1010
rect 12488 1178 12554 1194
rect 12488 1010 12504 1178
rect 12538 1010 12554 1178
rect 12488 960 12554 1010
rect 12608 1178 12674 1194
rect 12608 1010 12624 1178
rect 12658 1010 12674 1178
rect 12608 960 12674 1010
rect 12716 1178 12782 1430
rect 12818 1380 12884 1396
rect 12818 1346 12834 1380
rect 12868 1346 12884 1380
rect 12818 1330 12884 1346
rect 13052 1380 13118 1610
rect 13172 1678 13238 1728
rect 13172 1610 13188 1678
rect 13222 1610 13238 1678
rect 13172 1594 13238 1610
rect 13360 1678 13426 1694
rect 13360 1610 13376 1678
rect 13410 1610 13426 1678
rect 13360 1496 13426 1610
rect 13508 1678 13574 1728
rect 13508 1610 13524 1678
rect 13558 1610 13574 1678
rect 13508 1594 13574 1610
rect 13696 1678 13762 1694
rect 13696 1610 13712 1678
rect 13746 1610 13762 1678
rect 13696 1496 13762 1610
rect 13280 1430 13426 1496
rect 13616 1430 13762 1496
rect 13052 1346 13068 1380
rect 13102 1346 13118 1380
rect 13178 1410 13244 1426
rect 13178 1376 13194 1410
rect 13228 1376 13244 1410
rect 13178 1360 13244 1376
rect 13280 1410 13346 1430
rect 13280 1376 13296 1410
rect 13330 1376 13346 1410
rect 12950 1280 13016 1296
rect 12950 1246 12966 1280
rect 13000 1246 13016 1280
rect 12950 1230 13016 1246
rect 12716 1010 12732 1178
rect 12766 1010 12782 1178
rect 12716 994 12782 1010
rect 12824 1178 12890 1194
rect 12824 1010 12840 1178
rect 12874 1010 12890 1178
rect 12824 960 12890 1010
rect 12944 1178 13010 1194
rect 12944 1010 12960 1178
rect 12994 1010 13010 1178
rect 12944 960 13010 1010
rect 13052 1178 13118 1346
rect 13052 1010 13068 1178
rect 13102 1010 13118 1178
rect 13052 994 13118 1010
rect 13172 1178 13238 1194
rect 13172 1010 13188 1178
rect 13222 1010 13238 1178
rect 13172 960 13238 1010
rect 13280 1178 13346 1376
rect 13514 1410 13580 1426
rect 13514 1376 13530 1410
rect 13564 1376 13580 1410
rect 13514 1360 13580 1376
rect 13382 1328 13448 1344
rect 13382 1294 13398 1328
rect 13432 1294 13448 1328
rect 13382 1278 13448 1294
rect 13616 1328 13682 1430
rect 13616 1294 13632 1328
rect 13666 1294 13682 1328
rect 13280 1010 13296 1178
rect 13330 1010 13346 1178
rect 13280 994 13346 1010
rect 13388 1178 13454 1194
rect 13388 1010 13404 1178
rect 13438 1010 13454 1178
rect 13388 960 13454 1010
rect 13508 1178 13574 1194
rect 13508 1010 13524 1178
rect 13558 1010 13574 1178
rect 13508 960 13574 1010
rect 13616 1178 13682 1294
rect 13718 1328 13784 1344
rect 13718 1294 13734 1328
rect 13768 1294 13784 1328
rect 13718 1278 13784 1294
rect 13616 1010 13632 1178
rect 13666 1010 13682 1178
rect 13616 994 13682 1010
rect 13724 1178 13790 1194
rect 13724 1010 13740 1178
rect 13774 1010 13790 1178
rect 13724 960 13790 1010
rect 4 940 13862 960
rect 4 884 60 940
rect 266 884 368 940
rect 1838 884 1940 940
rect 3410 884 3512 940
rect 3718 884 3820 940
rect 5290 884 5392 940
rect 6862 884 6964 940
rect 7170 884 7272 940
rect 8742 884 8844 940
rect 10314 884 10416 940
rect 10622 884 10724 940
rect 12194 884 12296 940
rect 13766 884 13862 940
rect 4 864 13862 884
<< viali >>
rect 206 1493 250 1559
rect 884 1546 918 1580
rect 82 1410 148 1426
rect 82 1376 98 1410
rect 98 1376 132 1410
rect 132 1376 148 1410
rect 82 1360 148 1376
rect 614 1446 648 1480
rect 366 1246 400 1280
rect 641 1346 668 1375
rect 668 1346 675 1375
rect 641 1341 675 1346
rect 906 1346 940 1380
rect 1432 1563 1498 1597
rect 2456 1546 2490 1580
rect 2186 1446 2220 1480
rect 1140 1346 1174 1380
rect 1266 1376 1300 1410
rect 1368 1376 1402 1410
rect 1038 1246 1072 1280
rect 1602 1376 1636 1410
rect 1470 1294 1504 1328
rect 1704 1294 1738 1328
rect 1806 1294 1840 1328
rect 1938 1246 1972 1280
rect 2209 1380 2243 1381
rect 2209 1347 2240 1380
rect 2240 1347 2243 1380
rect 2478 1346 2512 1380
rect 3658 1493 3702 1559
rect 4336 1546 4370 1580
rect 2712 1346 2746 1380
rect 2838 1376 2872 1410
rect 2940 1376 2974 1410
rect 2610 1246 2644 1280
rect 3174 1376 3208 1410
rect 3042 1294 3076 1328
rect 3534 1410 3600 1426
rect 3534 1376 3550 1410
rect 3550 1376 3584 1410
rect 3584 1376 3600 1410
rect 3534 1360 3600 1376
rect 3276 1294 3310 1328
rect 3378 1294 3412 1328
rect 4066 1446 4100 1480
rect 3818 1246 3852 1280
rect 4093 1346 4120 1375
rect 4120 1346 4127 1375
rect 4093 1341 4127 1346
rect 4358 1346 4392 1380
rect 4884 1563 4950 1597
rect 5908 1546 5942 1580
rect 5638 1446 5672 1480
rect 4592 1346 4626 1380
rect 4718 1376 4752 1410
rect 4820 1376 4854 1410
rect 4490 1246 4524 1280
rect 5054 1376 5088 1410
rect 4922 1294 4956 1328
rect 5156 1294 5190 1328
rect 5258 1294 5292 1328
rect 5390 1246 5424 1280
rect 5661 1380 5695 1381
rect 5661 1347 5692 1380
rect 5692 1347 5695 1380
rect 5930 1346 5964 1380
rect 7110 1493 7154 1559
rect 7788 1546 7822 1580
rect 6164 1346 6198 1380
rect 6290 1376 6324 1410
rect 6392 1376 6426 1410
rect 6062 1246 6096 1280
rect 6626 1376 6660 1410
rect 6494 1294 6528 1328
rect 6986 1410 7052 1426
rect 6986 1376 7002 1410
rect 7002 1376 7036 1410
rect 7036 1376 7052 1410
rect 6986 1360 7052 1376
rect 6728 1294 6762 1328
rect 6830 1294 6864 1328
rect 7518 1446 7552 1480
rect 7270 1246 7304 1280
rect 7545 1346 7572 1375
rect 7572 1346 7579 1375
rect 7545 1341 7579 1346
rect 7810 1346 7844 1380
rect 8336 1563 8402 1597
rect 9360 1546 9394 1580
rect 9090 1446 9124 1480
rect 8044 1346 8078 1380
rect 8170 1376 8204 1410
rect 8272 1376 8306 1410
rect 7942 1246 7976 1280
rect 8506 1376 8540 1410
rect 8374 1294 8408 1328
rect 8608 1294 8642 1328
rect 8710 1294 8744 1328
rect 8842 1246 8876 1280
rect 9113 1380 9147 1381
rect 9113 1347 9144 1380
rect 9144 1347 9147 1380
rect 9382 1346 9416 1380
rect 10562 1493 10606 1559
rect 11240 1546 11274 1580
rect 9616 1346 9650 1380
rect 9742 1376 9776 1410
rect 9844 1376 9878 1410
rect 9514 1246 9548 1280
rect 10078 1376 10112 1410
rect 9946 1294 9980 1328
rect 10438 1410 10504 1426
rect 10438 1376 10454 1410
rect 10454 1376 10488 1410
rect 10488 1376 10504 1410
rect 10438 1360 10504 1376
rect 10180 1294 10214 1328
rect 10282 1294 10316 1328
rect 10970 1446 11004 1480
rect 10722 1246 10756 1280
rect 10997 1346 11024 1375
rect 11024 1346 11031 1375
rect 10997 1341 11031 1346
rect 11262 1346 11296 1380
rect 11788 1563 11854 1597
rect 12812 1546 12846 1580
rect 12542 1446 12576 1480
rect 11496 1346 11530 1380
rect 11622 1376 11656 1410
rect 11724 1376 11758 1410
rect 11394 1246 11428 1280
rect 11958 1376 11992 1410
rect 11826 1294 11860 1328
rect 12060 1294 12094 1328
rect 12162 1294 12196 1328
rect 12294 1246 12328 1280
rect 12565 1380 12599 1381
rect 12565 1347 12596 1380
rect 12596 1347 12599 1380
rect 12834 1346 12868 1380
rect 13068 1346 13102 1380
rect 13194 1376 13228 1410
rect 13296 1376 13330 1410
rect 12966 1246 13000 1280
rect 13530 1376 13564 1410
rect 13398 1294 13432 1328
rect 13632 1294 13666 1328
rect 13734 1294 13768 1328
<< metal1 >>
rect 408 1698 448 1700
rect 3860 1698 3900 1700
rect 7312 1698 7352 1700
rect 10764 1698 10804 1700
rect 408 1661 2068 1698
rect 200 1559 256 1571
rect 200 1493 206 1559
rect 250 1546 256 1559
rect 408 1546 448 1661
rect 1420 1597 1510 1603
rect 250 1506 448 1546
rect 868 1580 934 1594
rect 868 1546 884 1580
rect 918 1576 934 1580
rect 918 1546 1360 1576
rect 1420 1563 1432 1597
rect 1498 1594 1510 1597
rect 1498 1566 1974 1594
rect 1498 1563 1510 1566
rect 1420 1557 1510 1563
rect 868 1534 934 1546
rect 250 1493 256 1506
rect 200 1481 256 1493
rect 598 1480 664 1496
rect 1332 1486 1360 1546
rect 598 1446 614 1480
rect 648 1448 1300 1480
rect 1332 1456 1840 1486
rect 648 1446 664 1448
rect 76 1426 154 1438
rect 598 1430 664 1446
rect 76 1360 82 1426
rect 148 1415 154 1426
rect 1250 1426 1300 1448
rect 148 1381 340 1415
rect 1250 1410 1316 1426
rect 148 1375 687 1381
rect 148 1370 641 1375
rect 148 1360 154 1370
rect 76 1348 154 1360
rect 295 1341 641 1370
rect 675 1341 687 1375
rect 295 1336 687 1341
rect 629 1335 687 1336
rect 890 1380 956 1396
rect 1124 1380 1190 1396
rect 890 1346 906 1380
rect 940 1346 1140 1380
rect 1174 1346 1190 1380
rect 1250 1376 1266 1410
rect 1300 1376 1316 1410
rect 1250 1360 1316 1376
rect 1352 1410 1418 1426
rect 1586 1410 1652 1426
rect 1352 1376 1368 1410
rect 1402 1376 1602 1410
rect 1636 1376 1652 1410
rect 1352 1360 1418 1376
rect 1586 1360 1652 1376
rect 890 1330 956 1346
rect 1124 1330 1190 1346
rect 1806 1344 1840 1456
rect 1454 1328 1520 1344
rect 1688 1328 1754 1344
rect 350 1280 416 1296
rect 350 1246 366 1280
rect 400 1260 416 1280
rect 1022 1280 1088 1296
rect 1022 1260 1038 1280
rect 400 1246 1038 1260
rect 1072 1246 1088 1280
rect 1454 1294 1470 1328
rect 1504 1294 1704 1328
rect 1738 1294 1754 1328
rect 1454 1278 1520 1294
rect 1688 1278 1754 1294
rect 1790 1328 1856 1344
rect 1790 1294 1806 1328
rect 1840 1294 1856 1328
rect 1946 1296 1974 1566
rect 2031 1383 2068 1661
rect 3860 1661 5520 1698
rect 2440 1580 2506 1594
rect 2440 1546 2456 1580
rect 2490 1576 2506 1580
rect 2490 1546 2932 1576
rect 2440 1534 2506 1546
rect 2170 1480 2236 1496
rect 2904 1486 2932 1546
rect 3652 1559 3708 1571
rect 3652 1493 3658 1559
rect 3702 1546 3708 1559
rect 3860 1546 3900 1661
rect 4872 1597 4962 1603
rect 3702 1506 3900 1546
rect 4320 1580 4386 1594
rect 4320 1546 4336 1580
rect 4370 1576 4386 1580
rect 4370 1546 4812 1576
rect 4872 1563 4884 1597
rect 4950 1594 4962 1597
rect 4950 1566 5426 1594
rect 4950 1563 4962 1566
rect 4872 1557 4962 1563
rect 4320 1534 4386 1546
rect 3702 1493 3708 1506
rect 2170 1446 2186 1480
rect 2220 1448 2872 1480
rect 2904 1456 3412 1486
rect 3652 1481 3708 1493
rect 2220 1446 2236 1448
rect 2170 1430 2236 1446
rect 2822 1426 2872 1448
rect 2822 1410 2888 1426
rect 2197 1383 2255 1387
rect 2031 1381 2255 1383
rect 2031 1347 2209 1381
rect 2243 1347 2255 1381
rect 2031 1346 2255 1347
rect 2197 1341 2255 1346
rect 2462 1380 2528 1396
rect 2696 1380 2762 1396
rect 2462 1346 2478 1380
rect 2512 1346 2712 1380
rect 2746 1346 2762 1380
rect 2822 1376 2838 1410
rect 2872 1376 2888 1410
rect 2822 1360 2888 1376
rect 2924 1410 2990 1426
rect 3158 1410 3224 1426
rect 2924 1376 2940 1410
rect 2974 1376 3174 1410
rect 3208 1376 3224 1410
rect 2924 1360 2990 1376
rect 3158 1360 3224 1376
rect 2462 1330 2528 1346
rect 2696 1330 2762 1346
rect 3378 1344 3412 1456
rect 4050 1480 4116 1496
rect 4784 1486 4812 1546
rect 4050 1446 4066 1480
rect 4100 1448 4752 1480
rect 4784 1456 5292 1486
rect 4100 1446 4116 1448
rect 3528 1426 3606 1438
rect 4050 1430 4116 1446
rect 3528 1360 3534 1426
rect 3600 1415 3606 1426
rect 4702 1426 4752 1448
rect 3600 1381 3792 1415
rect 4702 1410 4768 1426
rect 3600 1375 4139 1381
rect 3600 1370 4093 1375
rect 3600 1360 3606 1370
rect 3528 1348 3606 1360
rect 3026 1328 3092 1344
rect 3260 1328 3326 1344
rect 1790 1278 1856 1294
rect 1922 1280 1988 1296
rect 350 1230 1088 1246
rect 1922 1246 1938 1280
rect 1972 1260 1988 1280
rect 2594 1280 2660 1296
rect 2594 1260 2610 1280
rect 1972 1246 2610 1260
rect 2644 1246 2660 1280
rect 3026 1294 3042 1328
rect 3076 1294 3276 1328
rect 3310 1294 3326 1328
rect 3026 1278 3092 1294
rect 3260 1278 3326 1294
rect 3362 1328 3428 1344
rect 3747 1341 4093 1370
rect 4127 1341 4139 1375
rect 3747 1336 4139 1341
rect 4081 1335 4139 1336
rect 4342 1380 4408 1396
rect 4576 1380 4642 1396
rect 4342 1346 4358 1380
rect 4392 1346 4592 1380
rect 4626 1346 4642 1380
rect 4702 1376 4718 1410
rect 4752 1376 4768 1410
rect 4702 1360 4768 1376
rect 4804 1410 4870 1426
rect 5038 1410 5104 1426
rect 4804 1376 4820 1410
rect 4854 1376 5054 1410
rect 5088 1376 5104 1410
rect 4804 1360 4870 1376
rect 5038 1360 5104 1376
rect 4342 1330 4408 1346
rect 4576 1330 4642 1346
rect 5258 1344 5292 1456
rect 3362 1294 3378 1328
rect 3412 1294 3428 1328
rect 4906 1328 4972 1344
rect 5140 1328 5206 1344
rect 3362 1278 3428 1294
rect 3802 1280 3868 1296
rect 1922 1230 2660 1246
rect 3802 1246 3818 1280
rect 3852 1260 3868 1280
rect 4474 1280 4540 1296
rect 4474 1260 4490 1280
rect 3852 1246 4490 1260
rect 4524 1246 4540 1280
rect 4906 1294 4922 1328
rect 4956 1294 5156 1328
rect 5190 1294 5206 1328
rect 4906 1278 4972 1294
rect 5140 1278 5206 1294
rect 5242 1328 5308 1344
rect 5242 1294 5258 1328
rect 5292 1294 5308 1328
rect 5398 1296 5426 1566
rect 5483 1383 5520 1661
rect 7312 1661 8972 1698
rect 5892 1580 5958 1594
rect 5892 1546 5908 1580
rect 5942 1576 5958 1580
rect 5942 1546 6384 1576
rect 5892 1534 5958 1546
rect 5622 1480 5688 1496
rect 6356 1486 6384 1546
rect 7104 1559 7160 1571
rect 7104 1493 7110 1559
rect 7154 1546 7160 1559
rect 7312 1546 7352 1661
rect 8324 1597 8414 1603
rect 7154 1506 7352 1546
rect 7772 1580 7838 1594
rect 7772 1546 7788 1580
rect 7822 1576 7838 1580
rect 7822 1546 8264 1576
rect 8324 1563 8336 1597
rect 8402 1594 8414 1597
rect 8402 1566 8878 1594
rect 8402 1563 8414 1566
rect 8324 1557 8414 1563
rect 7772 1534 7838 1546
rect 7154 1493 7160 1506
rect 5622 1446 5638 1480
rect 5672 1448 6324 1480
rect 6356 1456 6864 1486
rect 7104 1481 7160 1493
rect 5672 1446 5688 1448
rect 5622 1430 5688 1446
rect 6274 1426 6324 1448
rect 6274 1410 6340 1426
rect 5649 1383 5707 1387
rect 5483 1381 5707 1383
rect 5483 1347 5661 1381
rect 5695 1347 5707 1381
rect 5483 1346 5707 1347
rect 5649 1341 5707 1346
rect 5914 1380 5980 1396
rect 6148 1380 6214 1396
rect 5914 1346 5930 1380
rect 5964 1346 6164 1380
rect 6198 1346 6214 1380
rect 6274 1376 6290 1410
rect 6324 1376 6340 1410
rect 6274 1360 6340 1376
rect 6376 1410 6442 1426
rect 6610 1410 6676 1426
rect 6376 1376 6392 1410
rect 6426 1376 6626 1410
rect 6660 1376 6676 1410
rect 6376 1360 6442 1376
rect 6610 1360 6676 1376
rect 5914 1330 5980 1346
rect 6148 1330 6214 1346
rect 6830 1344 6864 1456
rect 7502 1480 7568 1496
rect 8236 1486 8264 1546
rect 7502 1446 7518 1480
rect 7552 1448 8204 1480
rect 8236 1456 8744 1486
rect 7552 1446 7568 1448
rect 6980 1426 7058 1438
rect 7502 1430 7568 1446
rect 6980 1360 6986 1426
rect 7052 1415 7058 1426
rect 8154 1426 8204 1448
rect 7052 1381 7244 1415
rect 8154 1410 8220 1426
rect 7052 1375 7591 1381
rect 7052 1370 7545 1375
rect 7052 1360 7058 1370
rect 6980 1348 7058 1360
rect 6478 1328 6544 1344
rect 6712 1328 6778 1344
rect 5242 1278 5308 1294
rect 5374 1280 5440 1296
rect 3802 1230 4540 1246
rect 5374 1246 5390 1280
rect 5424 1260 5440 1280
rect 6046 1280 6112 1296
rect 6046 1260 6062 1280
rect 5424 1246 6062 1260
rect 6096 1246 6112 1280
rect 6478 1294 6494 1328
rect 6528 1294 6728 1328
rect 6762 1294 6778 1328
rect 6478 1278 6544 1294
rect 6712 1278 6778 1294
rect 6814 1328 6880 1344
rect 7199 1341 7545 1370
rect 7579 1341 7591 1375
rect 7199 1336 7591 1341
rect 7533 1335 7591 1336
rect 7794 1380 7860 1396
rect 8028 1380 8094 1396
rect 7794 1346 7810 1380
rect 7844 1346 8044 1380
rect 8078 1346 8094 1380
rect 8154 1376 8170 1410
rect 8204 1376 8220 1410
rect 8154 1360 8220 1376
rect 8256 1410 8322 1426
rect 8490 1410 8556 1426
rect 8256 1376 8272 1410
rect 8306 1376 8506 1410
rect 8540 1376 8556 1410
rect 8256 1360 8322 1376
rect 8490 1360 8556 1376
rect 7794 1330 7860 1346
rect 8028 1330 8094 1346
rect 8710 1344 8744 1456
rect 6814 1294 6830 1328
rect 6864 1294 6880 1328
rect 8358 1328 8424 1344
rect 8592 1328 8658 1344
rect 6814 1278 6880 1294
rect 7254 1280 7320 1296
rect 5374 1230 6112 1246
rect 7254 1246 7270 1280
rect 7304 1260 7320 1280
rect 7926 1280 7992 1296
rect 7926 1260 7942 1280
rect 7304 1246 7942 1260
rect 7976 1246 7992 1280
rect 8358 1294 8374 1328
rect 8408 1294 8608 1328
rect 8642 1294 8658 1328
rect 8358 1278 8424 1294
rect 8592 1278 8658 1294
rect 8694 1328 8760 1344
rect 8694 1294 8710 1328
rect 8744 1294 8760 1328
rect 8850 1296 8878 1566
rect 8935 1383 8972 1661
rect 10764 1661 12424 1698
rect 9344 1580 9410 1594
rect 9344 1546 9360 1580
rect 9394 1576 9410 1580
rect 9394 1546 9836 1576
rect 9344 1534 9410 1546
rect 9074 1480 9140 1496
rect 9808 1486 9836 1546
rect 10556 1559 10612 1571
rect 10556 1493 10562 1559
rect 10606 1546 10612 1559
rect 10764 1546 10804 1661
rect 11776 1597 11866 1603
rect 10606 1506 10804 1546
rect 11224 1580 11290 1594
rect 11224 1546 11240 1580
rect 11274 1576 11290 1580
rect 11274 1546 11716 1576
rect 11776 1563 11788 1597
rect 11854 1594 11866 1597
rect 11854 1566 12330 1594
rect 11854 1563 11866 1566
rect 11776 1557 11866 1563
rect 11224 1534 11290 1546
rect 10606 1493 10612 1506
rect 9074 1446 9090 1480
rect 9124 1448 9776 1480
rect 9808 1456 10316 1486
rect 10556 1481 10612 1493
rect 9124 1446 9140 1448
rect 9074 1430 9140 1446
rect 9726 1426 9776 1448
rect 9726 1410 9792 1426
rect 9101 1383 9159 1387
rect 8935 1381 9159 1383
rect 8935 1347 9113 1381
rect 9147 1347 9159 1381
rect 8935 1346 9159 1347
rect 9101 1341 9159 1346
rect 9366 1380 9432 1396
rect 9600 1380 9666 1396
rect 9366 1346 9382 1380
rect 9416 1346 9616 1380
rect 9650 1346 9666 1380
rect 9726 1376 9742 1410
rect 9776 1376 9792 1410
rect 9726 1360 9792 1376
rect 9828 1410 9894 1426
rect 10062 1410 10128 1426
rect 9828 1376 9844 1410
rect 9878 1376 10078 1410
rect 10112 1376 10128 1410
rect 9828 1360 9894 1376
rect 10062 1360 10128 1376
rect 9366 1330 9432 1346
rect 9600 1330 9666 1346
rect 10282 1344 10316 1456
rect 10954 1480 11020 1496
rect 11688 1486 11716 1546
rect 10954 1446 10970 1480
rect 11004 1448 11656 1480
rect 11688 1456 12196 1486
rect 11004 1446 11020 1448
rect 10432 1426 10510 1438
rect 10954 1430 11020 1446
rect 10432 1360 10438 1426
rect 10504 1415 10510 1426
rect 11606 1426 11656 1448
rect 10504 1381 10696 1415
rect 11606 1410 11672 1426
rect 10504 1375 11043 1381
rect 10504 1370 10997 1375
rect 10504 1360 10510 1370
rect 10432 1348 10510 1360
rect 9930 1328 9996 1344
rect 10164 1328 10230 1344
rect 8694 1278 8760 1294
rect 8826 1280 8892 1296
rect 7254 1230 7992 1246
rect 8826 1246 8842 1280
rect 8876 1260 8892 1280
rect 9498 1280 9564 1296
rect 9498 1260 9514 1280
rect 8876 1246 9514 1260
rect 9548 1246 9564 1280
rect 9930 1294 9946 1328
rect 9980 1294 10180 1328
rect 10214 1294 10230 1328
rect 9930 1278 9996 1294
rect 10164 1278 10230 1294
rect 10266 1328 10332 1344
rect 10651 1341 10997 1370
rect 11031 1341 11043 1375
rect 10651 1336 11043 1341
rect 10985 1335 11043 1336
rect 11246 1380 11312 1396
rect 11480 1380 11546 1396
rect 11246 1346 11262 1380
rect 11296 1346 11496 1380
rect 11530 1346 11546 1380
rect 11606 1376 11622 1410
rect 11656 1376 11672 1410
rect 11606 1360 11672 1376
rect 11708 1410 11774 1426
rect 11942 1410 12008 1426
rect 11708 1376 11724 1410
rect 11758 1376 11958 1410
rect 11992 1376 12008 1410
rect 11708 1360 11774 1376
rect 11942 1360 12008 1376
rect 11246 1330 11312 1346
rect 11480 1330 11546 1346
rect 12162 1344 12196 1456
rect 10266 1294 10282 1328
rect 10316 1294 10332 1328
rect 11810 1328 11876 1344
rect 12044 1328 12110 1344
rect 10266 1278 10332 1294
rect 10706 1280 10772 1296
rect 8826 1230 9564 1246
rect 10706 1246 10722 1280
rect 10756 1260 10772 1280
rect 11378 1280 11444 1296
rect 11378 1260 11394 1280
rect 10756 1246 11394 1260
rect 11428 1246 11444 1280
rect 11810 1294 11826 1328
rect 11860 1294 12060 1328
rect 12094 1294 12110 1328
rect 11810 1278 11876 1294
rect 12044 1278 12110 1294
rect 12146 1328 12212 1344
rect 12146 1294 12162 1328
rect 12196 1294 12212 1328
rect 12302 1296 12330 1566
rect 12387 1383 12424 1661
rect 12796 1580 12862 1594
rect 12796 1546 12812 1580
rect 12846 1576 12862 1580
rect 12846 1546 13288 1576
rect 12796 1534 12862 1546
rect 12526 1480 12592 1496
rect 13260 1486 13288 1546
rect 12526 1446 12542 1480
rect 12576 1448 13228 1480
rect 13260 1456 13768 1486
rect 12576 1446 12592 1448
rect 12526 1430 12592 1446
rect 13178 1426 13228 1448
rect 13178 1410 13244 1426
rect 12553 1383 12611 1387
rect 12387 1381 12611 1383
rect 12387 1347 12565 1381
rect 12599 1347 12611 1381
rect 12387 1346 12611 1347
rect 12553 1341 12611 1346
rect 12818 1380 12884 1396
rect 13052 1380 13118 1396
rect 12818 1346 12834 1380
rect 12868 1346 13068 1380
rect 13102 1346 13118 1380
rect 13178 1376 13194 1410
rect 13228 1376 13244 1410
rect 13178 1360 13244 1376
rect 13280 1410 13346 1426
rect 13514 1410 13580 1426
rect 13280 1376 13296 1410
rect 13330 1376 13530 1410
rect 13564 1376 13580 1410
rect 13280 1360 13346 1376
rect 13514 1360 13580 1376
rect 12818 1330 12884 1346
rect 13052 1330 13118 1346
rect 13734 1344 13768 1456
rect 13382 1328 13448 1344
rect 13616 1328 13682 1344
rect 12146 1278 12212 1294
rect 12278 1280 12344 1296
rect 10706 1230 11444 1246
rect 12278 1246 12294 1280
rect 12328 1260 12344 1280
rect 12950 1280 13016 1296
rect 12950 1260 12966 1280
rect 12328 1246 12966 1260
rect 13000 1246 13016 1280
rect 13382 1294 13398 1328
rect 13432 1294 13632 1328
rect 13666 1294 13682 1328
rect 13382 1278 13448 1294
rect 13616 1278 13682 1294
rect 13718 1328 13784 1344
rect 13718 1294 13734 1328
rect 13768 1294 13784 1328
rect 13718 1278 13784 1294
rect 12278 1230 13016 1246
use DFF  DFF_0
timestamp 1681152781
transform 1 0 268 0 1 0
box -268 0 3242 976
use DFF  DFF_1
timestamp 1681152781
transform 1 0 3720 0 1 0
box -268 0 3242 976
use DFF  DFF_2
timestamp 1681152781
transform 1 0 7172 0 1 0
box -268 0 3242 976
use DFF  DFF_3
timestamp 1681152781
transform 1 0 10624 0 1 0
box -268 0 3242 976
<< labels >>
flabel locali s 10438 1360 10504 1426 0 FreeSerif 400 0 0 0 CLK
port 5 nsew
flabel locali 10360 1728 10678 1824 5 FreeSerif 160 0 0 0 GND!
port 1 n
flabel locali 10540 1194 10606 1594 5 FreeSerif 160 0 0 0 Y
port 2 n
flabel viali 10438 1360 10504 1426 0 FreeSerif 160 0 0 0 A
port 3 nsew
flabel locali 10360 864 10678 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali 12200 1728 13862 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 12200 864 13862 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 12278 1230 12344 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 12482 1330 12680 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 13360 1430 13426 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 13696 1430 13762 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 12344 1652 12344 1652 0 S$
rlabel ndiff 12424 1652 12424 1652 0 S$
rlabel ndiff 12680 1652 12680 1652 0 S$
rlabel ndiff 12760 1652 12760 1652 0 S$
rlabel ndiff 13016 1652 13016 1652 0 S$
rlabel ndiff 13244 1656 13244 1656 0 S$
rlabel ndiff 13324 1656 13324 1656 0 S$
rlabel ndiff 13580 1660 13580 1660 0 S$
rlabel ndiff 13660 1664 13660 1664 0 S$
rlabel pdiff 13718 1076 13718 1076 0 S$
rlabel pdiff 13580 1080 13580 1080 0 S$
rlabel pdiff 13382 1072 13382 1072 0 S$
rlabel pdiff 13244 1076 13244 1076 0 S$
rlabel pdiff 13016 1064 13016 1064 0 S$
rlabel pdiff 12818 1072 12818 1072 0 S$
rlabel pdiff 12680 1060 12680 1060 0 S$
rlabel pdiff 12482 1076 12482 1076 0 S$
rlabel pdiff 12344 1072 12344 1072 0 S$
flabel locali 10628 1728 12290 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 10628 864 12290 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 10706 1230 10772 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 10910 1330 11108 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 11788 1430 11854 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 12124 1430 12190 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 10772 1652 10772 1652 0 S$
rlabel ndiff 10852 1652 10852 1652 0 S$
rlabel ndiff 11108 1652 11108 1652 0 S$
rlabel ndiff 11188 1652 11188 1652 0 S$
rlabel ndiff 11444 1652 11444 1652 0 S$
rlabel ndiff 11672 1656 11672 1656 0 S$
rlabel ndiff 11752 1656 11752 1656 0 S$
rlabel ndiff 12008 1660 12008 1660 0 S$
rlabel ndiff 12088 1664 12088 1664 0 S$
rlabel pdiff 12146 1076 12146 1076 0 S$
rlabel pdiff 12008 1080 12008 1080 0 S$
rlabel pdiff 11810 1072 11810 1072 0 S$
rlabel pdiff 11672 1076 11672 1076 0 S$
rlabel pdiff 11444 1064 11444 1064 0 S$
rlabel pdiff 11246 1072 11246 1072 0 S$
rlabel pdiff 11108 1060 11108 1060 0 S$
rlabel pdiff 10910 1076 10910 1076 0 S$
rlabel pdiff 10772 1072 10772 1072 0 S$
flabel locali s 6986 1360 7052 1426 0 FreeSerif 400 0 0 0 CLK
port 5 nsew
flabel locali 6908 1728 7226 1824 5 FreeSerif 160 0 0 0 GND!
port 1 n
flabel locali 7088 1194 7154 1594 5 FreeSerif 160 0 0 0 Y
port 2 n
flabel viali 6986 1360 7052 1426 0 FreeSerif 160 0 0 0 A
port 3 nsew
flabel locali 6908 864 7226 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali 8748 1728 10410 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 8748 864 10410 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 8826 1230 8892 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 9030 1330 9228 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 9908 1430 9974 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 10244 1430 10310 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 8892 1652 8892 1652 0 S$
rlabel ndiff 8972 1652 8972 1652 0 S$
rlabel ndiff 9228 1652 9228 1652 0 S$
rlabel ndiff 9308 1652 9308 1652 0 S$
rlabel ndiff 9564 1652 9564 1652 0 S$
rlabel ndiff 9792 1656 9792 1656 0 S$
rlabel ndiff 9872 1656 9872 1656 0 S$
rlabel ndiff 10128 1660 10128 1660 0 S$
rlabel ndiff 10208 1664 10208 1664 0 S$
rlabel pdiff 10266 1076 10266 1076 0 S$
rlabel pdiff 10128 1080 10128 1080 0 S$
rlabel pdiff 9930 1072 9930 1072 0 S$
rlabel pdiff 9792 1076 9792 1076 0 S$
rlabel pdiff 9564 1064 9564 1064 0 S$
rlabel pdiff 9366 1072 9366 1072 0 S$
rlabel pdiff 9228 1060 9228 1060 0 S$
rlabel pdiff 9030 1076 9030 1076 0 S$
rlabel pdiff 8892 1072 8892 1072 0 S$
flabel locali 7176 1728 8838 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 7176 864 8838 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 7254 1230 7320 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 7458 1330 7656 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 8336 1430 8402 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 8672 1430 8738 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 7320 1652 7320 1652 0 S$
rlabel ndiff 7400 1652 7400 1652 0 S$
rlabel ndiff 7656 1652 7656 1652 0 S$
rlabel ndiff 7736 1652 7736 1652 0 S$
rlabel ndiff 7992 1652 7992 1652 0 S$
rlabel ndiff 8220 1656 8220 1656 0 S$
rlabel ndiff 8300 1656 8300 1656 0 S$
rlabel ndiff 8556 1660 8556 1660 0 S$
rlabel ndiff 8636 1664 8636 1664 0 S$
rlabel pdiff 8694 1076 8694 1076 0 S$
rlabel pdiff 8556 1080 8556 1080 0 S$
rlabel pdiff 8358 1072 8358 1072 0 S$
rlabel pdiff 8220 1076 8220 1076 0 S$
rlabel pdiff 7992 1064 7992 1064 0 S$
rlabel pdiff 7794 1072 7794 1072 0 S$
rlabel pdiff 7656 1060 7656 1060 0 S$
rlabel pdiff 7458 1076 7458 1076 0 S$
rlabel pdiff 7320 1072 7320 1072 0 S$
flabel locali s 3534 1360 3600 1426 0 FreeSerif 400 0 0 0 CLK
port 5 nsew
flabel locali 3456 1728 3774 1824 5 FreeSerif 160 0 0 0 GND!
port 1 n
flabel locali 3636 1194 3702 1594 5 FreeSerif 160 0 0 0 Y
port 2 n
flabel viali 3534 1360 3600 1426 0 FreeSerif 160 0 0 0 A
port 3 nsew
flabel locali 3456 864 3774 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali 5296 1728 6958 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 5296 864 6958 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 5374 1230 5440 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 5578 1330 5776 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 6456 1430 6522 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 6792 1430 6858 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 5440 1652 5440 1652 0 S$
rlabel ndiff 5520 1652 5520 1652 0 S$
rlabel ndiff 5776 1652 5776 1652 0 S$
rlabel ndiff 5856 1652 5856 1652 0 S$
rlabel ndiff 6112 1652 6112 1652 0 S$
rlabel ndiff 6340 1656 6340 1656 0 S$
rlabel ndiff 6420 1656 6420 1656 0 S$
rlabel ndiff 6676 1660 6676 1660 0 S$
rlabel ndiff 6756 1664 6756 1664 0 S$
rlabel pdiff 6814 1076 6814 1076 0 S$
rlabel pdiff 6676 1080 6676 1080 0 S$
rlabel pdiff 6478 1072 6478 1072 0 S$
rlabel pdiff 6340 1076 6340 1076 0 S$
rlabel pdiff 6112 1064 6112 1064 0 S$
rlabel pdiff 5914 1072 5914 1072 0 S$
rlabel pdiff 5776 1060 5776 1060 0 S$
rlabel pdiff 5578 1076 5578 1076 0 S$
rlabel pdiff 5440 1072 5440 1072 0 S$
flabel locali 3724 1728 5386 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 3724 864 5386 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 3802 1230 3868 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 4006 1330 4204 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 4884 1430 4950 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 5220 1430 5286 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 3868 1652 3868 1652 0 S$
rlabel ndiff 3948 1652 3948 1652 0 S$
rlabel ndiff 4204 1652 4204 1652 0 S$
rlabel ndiff 4284 1652 4284 1652 0 S$
rlabel ndiff 4540 1652 4540 1652 0 S$
rlabel ndiff 4768 1656 4768 1656 0 S$
rlabel ndiff 4848 1656 4848 1656 0 S$
rlabel ndiff 5104 1660 5104 1660 0 S$
rlabel ndiff 5184 1664 5184 1664 0 S$
rlabel pdiff 5242 1076 5242 1076 0 S$
rlabel pdiff 5104 1080 5104 1080 0 S$
rlabel pdiff 4906 1072 4906 1072 0 S$
rlabel pdiff 4768 1076 4768 1076 0 S$
rlabel pdiff 4540 1064 4540 1064 0 S$
rlabel pdiff 4342 1072 4342 1072 0 S$
rlabel pdiff 4204 1060 4204 1060 0 S$
rlabel pdiff 4006 1076 4006 1076 0 S$
rlabel pdiff 3868 1072 3868 1072 0 S$
flabel locali s 82 1360 148 1426 0 FreeSerif 400 0 0 0 CLK
port 5 nsew
flabel locali 4 1728 322 1824 5 FreeSerif 160 0 0 0 GND!
port 1 n
flabel locali 184 1194 250 1594 5 FreeSerif 160 0 0 0 Y
port 2 n
flabel viali 82 1360 148 1426 0 FreeSerif 160 0 0 0 A
port 3 nsew
flabel locali 4 864 322 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali 1844 1728 3506 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 1844 864 3506 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 1922 1230 1988 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 2126 1330 2324 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 3004 1430 3070 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 3340 1430 3406 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 1988 1652 1988 1652 0 S$
rlabel ndiff 2068 1652 2068 1652 0 S$
rlabel ndiff 2324 1652 2324 1652 0 S$
rlabel ndiff 2404 1652 2404 1652 0 S$
rlabel ndiff 2660 1652 2660 1652 0 S$
rlabel ndiff 2888 1656 2888 1656 0 S$
rlabel ndiff 2968 1656 2968 1656 0 S$
rlabel ndiff 3224 1660 3224 1660 0 S$
rlabel ndiff 3304 1664 3304 1664 0 S$
rlabel pdiff 3362 1076 3362 1076 0 S$
rlabel pdiff 3224 1080 3224 1080 0 S$
rlabel pdiff 3026 1072 3026 1072 0 S$
rlabel pdiff 2888 1076 2888 1076 0 S$
rlabel pdiff 2660 1064 2660 1064 0 S$
rlabel pdiff 2462 1072 2462 1072 0 S$
rlabel pdiff 2324 1060 2324 1060 0 S$
rlabel pdiff 2126 1076 2126 1076 0 S$
rlabel pdiff 1988 1072 1988 1072 0 S$
flabel locali 272 1728 1934 1824 0 FreeSerif 160 0 0 0 GND!
port 11 nsew
flabel locali 272 864 1934 960 0 FreeSerif 160 0 0 0 VDD!
port 0 nsew
flabel locali s 350 1230 416 1296 0 FreeSerif 160 0 0 0 D
port 1 nsew
flabel locali s 554 1330 752 1396 0 FreeSerif 160 0 0 0 CLK
port 6 nsew
flabel locali s 1432 1430 1498 1594 0 FreeSerif 160 0 0 0 Q
port 22 nsew
flabel locali s 1768 1430 1834 1594 0 FreeSerif 160 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 416 1652 416 1652 0 S$
rlabel ndiff 496 1652 496 1652 0 S$
rlabel ndiff 752 1652 752 1652 0 S$
rlabel ndiff 832 1652 832 1652 0 S$
rlabel ndiff 1088 1652 1088 1652 0 S$
rlabel ndiff 1316 1656 1316 1656 0 S$
rlabel ndiff 1396 1656 1396 1656 0 S$
rlabel ndiff 1652 1660 1652 1660 0 S$
rlabel ndiff 1732 1664 1732 1664 0 S$
rlabel pdiff 1790 1076 1790 1076 0 S$
rlabel pdiff 1652 1080 1652 1080 0 S$
rlabel pdiff 1454 1072 1454 1072 0 S$
rlabel pdiff 1316 1076 1316 1076 0 S$
rlabel pdiff 1088 1064 1088 1064 0 S$
rlabel pdiff 890 1072 890 1072 0 S$
rlabel pdiff 752 1060 752 1060 0 S$
rlabel pdiff 554 1076 554 1076 0 S$
rlabel pdiff 416 1072 416 1072 0 S$
<< end >>
