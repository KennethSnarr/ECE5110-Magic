* NGSPICE file created from nand2.ext - technology: sky130A

*.subckt nand2 VDD GND Y A B
X0 a_94_6# A GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=7.2e+11p pd=5.44e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X2 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B a_94_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
*.ends

