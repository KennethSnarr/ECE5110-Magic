magic
tech sky130A
magscale 1 2
timestamp 1681434240
<< locali >>
rect -264 864 8158 960
rect -186 398 -120 423
rect -84 321 -18 630
rect 82 398 148 464
rect 184 449 250 630
rect 286 537 352 546
rect 286 503 305 537
rect 339 503 352 537
rect 286 480 352 503
rect 184 415 204 449
rect 238 415 250 449
rect 184 328 250 415
rect 453 398 484 464
rect 520 328 586 630
rect 622 480 654 546
rect 856 530 922 630
rect 856 496 869 530
rect 903 496 922 530
rect 754 447 820 464
rect 754 413 773 447
rect 807 413 820 447
rect 754 398 820 413
rect 856 328 922 496
rect 958 480 1024 546
rect 1090 398 1156 464
rect 1192 449 1258 630
rect 1294 532 1360 546
rect 1294 498 1307 532
rect 1341 498 1360 532
rect 1294 480 1360 498
rect 1192 415 1212 449
rect 1246 415 1258 449
rect 1192 328 1258 415
rect 1461 398 1492 464
rect 1528 328 1594 630
rect 1630 480 1662 546
rect 1864 530 1930 630
rect 1864 496 1877 530
rect 1911 496 1930 530
rect 1762 447 1828 464
rect 1762 413 1783 447
rect 1817 413 1828 447
rect 1762 398 1828 413
rect 1864 328 1930 496
rect 1966 480 2032 546
rect 2098 398 2164 464
rect 2200 449 2266 630
rect 2302 530 2368 546
rect 2302 496 2315 530
rect 2349 496 2368 530
rect 2302 480 2368 496
rect 2200 415 2220 449
rect 2254 415 2266 449
rect 2200 328 2266 415
rect 2469 398 2500 464
rect 2536 328 2602 630
rect 2638 480 2670 546
rect 2872 530 2938 630
rect 2872 496 2885 530
rect 2919 496 2938 530
rect 2770 449 2836 464
rect 2770 415 2787 449
rect 2821 415 2836 449
rect 2770 398 2836 415
rect 2872 328 2938 496
rect 2974 480 3040 546
rect 3106 398 3172 464
rect 3208 449 3274 630
rect 3310 532 3376 546
rect 3310 498 3319 532
rect 3353 498 3376 532
rect 3310 480 3376 498
rect 3208 415 3228 449
rect 3262 415 3274 449
rect 3208 328 3274 415
rect 3477 398 3508 464
rect 3544 328 3610 630
rect 3646 480 3678 546
rect 3880 530 3946 630
rect 3880 496 3893 530
rect 3927 496 3946 530
rect 3778 447 3844 464
rect 3778 413 3799 447
rect 3833 413 3844 447
rect 3778 398 3844 413
rect 3880 328 3946 496
rect 3982 480 4048 546
rect 4114 398 4180 464
rect 4216 449 4282 630
rect 4318 530 4384 546
rect 4318 496 4331 530
rect 4365 496 4384 530
rect 4318 480 4384 496
rect 4216 415 4236 449
rect 4270 415 4282 449
rect 4216 328 4282 415
rect 4485 398 4516 464
rect 4552 328 4618 630
rect 4654 480 4686 546
rect 4888 530 4954 630
rect 4888 496 4901 530
rect 4935 496 4954 530
rect 4786 449 4852 464
rect 4786 415 4807 449
rect 4841 415 4852 449
rect 4786 398 4852 415
rect 4888 328 4954 496
rect 4990 480 5056 546
rect 5122 398 5188 464
rect 5224 449 5290 630
rect 5326 528 5392 546
rect 5326 494 5341 528
rect 5375 494 5392 528
rect 5326 480 5392 494
rect 5224 415 5244 449
rect 5278 415 5290 449
rect 5224 328 5290 415
rect 5493 398 5524 464
rect 5560 328 5626 630
rect 5662 480 5694 546
rect 5896 530 5962 630
rect 5896 496 5909 530
rect 5943 496 5962 530
rect 5794 449 5860 464
rect 5794 415 5807 449
rect 5841 415 5860 449
rect 5794 398 5860 415
rect 5896 328 5962 496
rect 5998 480 6064 546
rect 6130 398 6196 464
rect 6232 449 6298 630
rect 6334 536 6400 546
rect 6334 502 6351 536
rect 6385 502 6400 536
rect 6334 480 6400 502
rect 6232 415 6252 449
rect 6286 415 6298 449
rect 6232 328 6298 415
rect 6501 398 6532 464
rect 6568 328 6634 630
rect 6670 480 6702 546
rect 6904 530 6970 630
rect 6904 496 6917 530
rect 6951 496 6970 530
rect 6802 447 6868 464
rect 6802 413 6821 447
rect 6855 413 6868 447
rect 6802 398 6868 413
rect 6904 328 6970 496
rect 7006 480 7072 546
rect 7138 398 7204 464
rect 7240 449 7306 630
rect 7342 538 7408 546
rect 7342 504 7357 538
rect 7391 504 7408 538
rect 7342 480 7408 504
rect 7240 415 7260 449
rect 7294 415 7306 449
rect 7240 328 7306 415
rect 7509 398 7540 464
rect 7576 328 7642 630
rect 7678 480 7710 546
rect 7912 530 7978 630
rect 7912 496 7925 530
rect 7959 496 7978 530
rect 7810 451 7876 464
rect 7810 417 7825 451
rect 7859 417 7876 451
rect 7810 398 7876 417
rect 7912 328 7978 496
rect 8014 480 8080 546
rect -84 255 -53 321
rect -84 230 -18 255
rect -264 0 8158 96
<< viali >>
rect -186 423 -120 464
rect 305 503 339 537
rect 204 415 238 449
rect 418 398 453 464
rect 654 480 688 546
rect 869 496 903 530
rect 773 413 807 447
rect 1307 498 1341 532
rect 1212 415 1246 449
rect 1426 398 1461 464
rect 1662 480 1696 546
rect 1877 496 1911 530
rect 1783 413 1817 447
rect 2315 496 2349 530
rect 2220 415 2254 449
rect 2434 398 2469 464
rect 2670 480 2704 546
rect 2885 496 2919 530
rect 2787 415 2821 449
rect 3319 498 3353 532
rect 3228 415 3262 449
rect 3442 398 3477 464
rect 3678 480 3712 546
rect 3893 496 3927 530
rect 3799 413 3833 447
rect 4331 496 4365 530
rect 4236 415 4270 449
rect 4450 398 4485 464
rect 4686 480 4720 546
rect 4901 496 4935 530
rect 4807 415 4841 449
rect 5341 494 5375 528
rect 5244 415 5278 449
rect 5458 398 5493 464
rect 5694 480 5728 546
rect 5909 496 5943 530
rect 5807 415 5841 449
rect 6351 502 6385 536
rect 6252 415 6286 449
rect 6466 398 6501 464
rect 6702 480 6736 546
rect 6917 496 6951 530
rect 6821 413 6855 447
rect 7357 504 7391 538
rect 7260 415 7294 449
rect 7474 398 7509 464
rect 7710 480 7744 546
rect 7925 496 7959 530
rect 7825 417 7859 451
rect -53 255 -18 321
<< metal1 >>
rect 305 589 7390 622
rect 305 543 338 589
rect 648 546 694 558
rect 293 537 351 543
rect 293 536 305 537
rect -169 503 305 536
rect 339 503 351 537
rect -169 470 -136 503
rect 293 497 351 503
rect 648 480 654 546
rect 688 530 694 546
rect 1307 544 1340 589
rect 1656 546 1702 558
rect 857 530 915 536
rect 688 496 869 530
rect 903 496 915 530
rect 688 480 694 496
rect 857 490 915 496
rect 1301 532 1347 544
rect 1301 498 1307 532
rect 1341 498 1347 532
rect 1301 486 1347 498
rect -198 464 -108 470
rect -198 423 -186 464
rect -120 423 -108 464
rect 412 464 459 476
rect 648 468 694 480
rect 1656 480 1662 546
rect 1696 530 1702 546
rect 2315 542 2348 589
rect 2664 546 2710 558
rect 1865 530 1923 536
rect 1696 496 1877 530
rect 1911 496 1923 530
rect 1696 480 1702 496
rect 1865 490 1923 496
rect 2309 530 2355 542
rect 2309 496 2315 530
rect 2349 496 2355 530
rect 2309 484 2355 496
rect -198 417 -108 423
rect 192 449 250 455
rect 412 449 418 464
rect 192 415 204 449
rect 238 415 418 449
rect 192 414 418 415
rect 192 409 250 414
rect 412 398 418 414
rect 453 398 459 464
rect 1420 464 1467 476
rect 1656 468 1702 480
rect 2664 480 2670 546
rect 2704 530 2710 546
rect 3319 544 3352 589
rect 3672 546 3718 558
rect 2873 530 2931 536
rect 2704 496 2885 530
rect 2919 496 2931 530
rect 2704 480 2710 496
rect 2873 490 2931 496
rect 3313 532 3359 544
rect 3313 498 3319 532
rect 3353 498 3359 532
rect 3313 486 3359 498
rect 767 447 813 459
rect 767 413 773 447
rect 807 413 813 447
rect 767 401 813 413
rect 1200 449 1258 455
rect 1420 449 1426 464
rect 1200 415 1212 449
rect 1246 415 1426 449
rect 1200 414 1426 415
rect 1200 409 1258 414
rect 412 386 459 398
rect -59 321 -12 333
rect -59 255 -53 321
rect -18 306 -12 321
rect 772 306 807 401
rect 1420 398 1426 414
rect 1461 398 1467 464
rect 2428 464 2475 476
rect 2664 468 2710 480
rect 3672 480 3678 546
rect 3712 530 3718 546
rect 4331 542 4364 589
rect 4680 546 4726 558
rect 3881 530 3939 536
rect 3712 496 3893 530
rect 3927 496 3939 530
rect 3712 480 3718 496
rect 3881 490 3939 496
rect 4325 530 4371 542
rect 4325 496 4331 530
rect 4365 496 4371 530
rect 4325 484 4371 496
rect 1777 447 1823 459
rect 1777 413 1783 447
rect 1817 413 1823 447
rect 1777 401 1823 413
rect 2208 449 2266 455
rect 2428 449 2434 464
rect 2208 415 2220 449
rect 2254 415 2434 449
rect 2208 414 2434 415
rect 2208 409 2266 414
rect 1420 386 1467 398
rect 1782 306 1817 401
rect 2428 398 2434 414
rect 2469 398 2475 464
rect 3436 464 3483 476
rect 3672 468 3718 480
rect 4680 480 4686 546
rect 4720 530 4726 546
rect 5341 540 5374 589
rect 5688 546 5734 558
rect 6351 548 6384 589
rect 4889 530 4947 536
rect 4720 496 4901 530
rect 4935 496 4947 530
rect 4720 480 4726 496
rect 4889 490 4947 496
rect 5335 528 5381 540
rect 5335 494 5341 528
rect 5375 494 5381 528
rect 5335 482 5381 494
rect 2781 449 2827 461
rect 2781 415 2787 449
rect 2821 415 2827 449
rect 2781 403 2827 415
rect 3216 449 3274 455
rect 3436 449 3442 464
rect 3216 415 3228 449
rect 3262 415 3442 449
rect 3216 414 3442 415
rect 3216 409 3274 414
rect 2428 386 2475 398
rect 2786 307 2821 403
rect 3436 398 3442 414
rect 3477 398 3483 464
rect 4444 464 4491 476
rect 4680 468 4726 480
rect 5688 480 5694 546
rect 5728 530 5734 546
rect 6345 536 6391 548
rect 5897 530 5955 536
rect 5728 496 5909 530
rect 5943 496 5955 530
rect 5728 480 5734 496
rect 5897 490 5955 496
rect 6345 502 6351 536
rect 6385 502 6391 536
rect 6345 490 6391 502
rect 6696 546 6742 558
rect 7357 550 7390 589
rect 3793 447 3839 459
rect 3793 413 3799 447
rect 3833 413 3839 447
rect 3793 401 3839 413
rect 4224 449 4282 455
rect 4444 449 4450 464
rect 4224 415 4236 449
rect 4270 415 4450 449
rect 4224 414 4450 415
rect 4224 409 4282 414
rect 3436 386 3483 398
rect 3798 307 3833 401
rect 4444 398 4450 414
rect 4485 398 4491 464
rect 5452 464 5499 476
rect 5688 468 5734 480
rect 6696 480 6702 546
rect 6736 530 6742 546
rect 7351 538 7397 550
rect 6905 530 6963 536
rect 6736 496 6917 530
rect 6951 496 6963 530
rect 6736 480 6742 496
rect 6905 490 6963 496
rect 7351 504 7357 538
rect 7391 504 7397 538
rect 7351 492 7397 504
rect 7704 546 7750 558
rect 4801 449 4847 461
rect 4801 415 4807 449
rect 4841 415 4847 449
rect 4801 403 4847 415
rect 5232 449 5290 455
rect 5452 449 5458 464
rect 5232 415 5244 449
rect 5278 415 5458 449
rect 5232 414 5458 415
rect 5232 409 5290 414
rect 4444 386 4491 398
rect 4806 307 4841 403
rect 5452 398 5458 414
rect 5493 398 5499 464
rect 6460 464 6507 476
rect 6696 468 6742 480
rect 7704 480 7710 546
rect 7744 530 7750 546
rect 7913 530 7971 536
rect 7744 496 7925 530
rect 7959 496 7971 530
rect 7744 480 7750 496
rect 7913 490 7971 496
rect 5801 449 5847 461
rect 5801 415 5807 449
rect 5841 415 5847 449
rect 5801 403 5847 415
rect 6240 449 6298 455
rect 6460 449 6466 464
rect 6240 415 6252 449
rect 6286 415 6466 449
rect 6240 414 6466 415
rect 6240 409 6298 414
rect 5452 386 5499 398
rect 5806 307 5841 403
rect 6460 398 6466 414
rect 6501 398 6507 464
rect 7468 464 7515 476
rect 7704 468 7750 480
rect 6815 447 6861 459
rect 6815 413 6821 447
rect 6855 413 6861 447
rect 6815 401 6861 413
rect 7248 449 7306 455
rect 7468 449 7474 464
rect 7248 415 7260 449
rect 7294 415 7474 449
rect 7248 414 7474 415
rect 7248 409 7306 414
rect 6460 386 6507 398
rect 6820 307 6855 401
rect 7468 398 7474 414
rect 7509 398 7515 464
rect 7819 451 7865 463
rect 7819 417 7825 451
rect 7859 417 7865 451
rect 7819 405 7865 417
rect 7468 386 7515 398
rect 7824 307 7859 405
rect 2786 306 7859 307
rect -18 272 7859 306
rect -18 271 2821 272
rect -18 255 -12 271
rect -59 243 -12 255
use inv  inv_0
timestamp 1679616770
transform 1 0 -184 0 1 124
box -84 -124 242 852
use nand2  nand2_0
timestamp 1676660346
transform 1 0 84 0 1 124
box -84 -124 350 852
use nand2  nand2_1
timestamp 1676660346
transform 1 0 420 0 1 124
box -84 -124 350 852
use nand2  nand2_2
timestamp 1676660346
transform 1 0 756 0 1 124
box -84 -124 350 852
use nand2  nand2_3
timestamp 1676660346
transform 1 0 1764 0 1 124
box -84 -124 350 852
use nand2  nand2_4
timestamp 1676660346
transform 1 0 1428 0 1 124
box -84 -124 350 852
use nand2  nand2_5
timestamp 1676660346
transform 1 0 1092 0 1 124
box -84 -124 350 852
use nand2  nand2_6
timestamp 1676660346
transform 1 0 2100 0 1 124
box -84 -124 350 852
use nand2  nand2_7
timestamp 1676660346
transform 1 0 2436 0 1 124
box -84 -124 350 852
use nand2  nand2_8
timestamp 1676660346
transform 1 0 2772 0 1 124
box -84 -124 350 852
use nand2  nand2_9
timestamp 1676660346
transform 1 0 3108 0 1 124
box -84 -124 350 852
use nand2  nand2_10
timestamp 1676660346
transform 1 0 3444 0 1 124
box -84 -124 350 852
use nand2  nand2_11
timestamp 1676660346
transform 1 0 3780 0 1 124
box -84 -124 350 852
use nand2  nand2_12
timestamp 1676660346
transform 1 0 4116 0 1 124
box -84 -124 350 852
use nand2  nand2_13
timestamp 1676660346
transform 1 0 4452 0 1 124
box -84 -124 350 852
use nand2  nand2_14
timestamp 1676660346
transform 1 0 4788 0 1 124
box -84 -124 350 852
use nand2  nand2_15
timestamp 1676660346
transform 1 0 5124 0 1 124
box -84 -124 350 852
use nand2  nand2_16
timestamp 1676660346
transform 1 0 5460 0 1 124
box -84 -124 350 852
use nand2  nand2_17
timestamp 1676660346
transform 1 0 5796 0 1 124
box -84 -124 350 852
use nand2  nand2_18
timestamp 1676660346
transform 1 0 6132 0 1 124
box -84 -124 350 852
use nand2  nand2_19
timestamp 1676660346
transform 1 0 6468 0 1 124
box -84 -124 350 852
use nand2  nand2_20
timestamp 1676660346
transform 1 0 7140 0 1 124
box -84 -124 350 852
use nand2  nand2_21
timestamp 1676660346
transform 1 0 6804 0 1 124
box -84 -124 350 852
use nand2  nand2_22
timestamp 1676660346
transform 1 0 7476 0 1 124
box -84 -124 350 852
use nand2  nand2_23
timestamp 1676660346
transform 1 0 7812 0 1 124
box -84 -124 350 852
<< labels >>
flabel locali s 520 328 586 630 0 FreeSerif 240 0 0 0 Y0
port 16 nsew
flabel locali s 82 398 148 464 0 FreeSerif 400 0 0 0 A0
port 15 nsew
flabel locali s 958 480 1024 546 0 FreeSerif 400 0 0 0 B0
port 17 nsew
flabel locali s 1090 398 1156 464 0 FreeSerif 400 0 0 0 A1
port 21 nsew
flabel locali s 1966 480 2032 546 0 FreeSerif 400 0 0 0 B1
port 23 nsew
flabel locali s 2098 398 2164 464 0 FreeSerif 400 0 0 0 A2
port 3 nsew
flabel locali s 2974 480 3040 546 0 FreeSerif 400 0 0 0 B2
port 5 nsew
flabel locali s 3106 398 3172 464 0 FreeSerif 400 0 0 0 A3
port 9 nsew
flabel locali s 3982 480 4048 546 0 FreeSerif 400 0 0 0 B3
port 11 nsew
flabel locali s 4114 398 4180 464 0 FreeSerif 400 0 0 0 A4
port 39 nsew
flabel locali s 4990 480 5056 546 0 FreeSerif 400 0 0 0 B4
port 41 nsew
flabel locali s 5122 398 5188 464 0 FreeSerif 400 0 0 0 A5
port 45 nsew
flabel locali s 5998 480 6064 546 0 FreeSerif 400 0 0 0 B5
port 47 nsew
flabel locali s 6130 398 6196 464 0 FreeSerif 400 0 0 0 A6
port 27 nsew
flabel locali s 7006 480 7072 546 0 FreeSerif 400 0 0 0 B6
port 29 nsew
flabel locali s 7138 398 7204 464 0 FreeSerif 400 0 0 0 A7
port 33 nsew
flabel locali s 8014 480 8080 546 0 FreeSerif 400 0 0 0 B7
port 35 nsew
flabel locali s -186 398 -120 464 0 FreeSerif 400 0 0 0 SEL
port 48 nsew
flabel locali s 1528 328 1594 630 0 FreeSerif 400 0 0 0 Y1
port 22 nsew
flabel locali s 2536 328 2602 630 0 FreeSerif 400 0 0 0 Y2
port 4 nsew
flabel locali s 3544 328 3610 630 0 FreeSerif 400 0 0 0 Y3
port 10 nsew
flabel locali s 4552 328 4618 630 0 FreeSerif 400 0 0 0 Y4
port 40 nsew
flabel locali s 5560 328 5626 630 0 FreeSerif 400 0 0 0 Y5
port 46 nsew
flabel locali s 6568 328 6634 630 0 FreeSerif 400 0 0 0 Y6
port 28 nsew
flabel locali s 7576 328 7642 630 0 FreeSerif 400 0 0 0 Y7
port 34 nsew
flabel locali s -264 864 8158 960 0 FreeSerif 400 0 0 0 VDD!
flabel locali s -264 0 8158 96 0 FreeSerif 400 0 0 0 GND!
<< end >>
