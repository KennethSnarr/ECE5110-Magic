* NGSPICE file created from multiplexor.ext - technology: sky130A

.subckt nand2 VDD GND Y A B
X0 a_94_6# A GND GND sky130_fd_pr__nfet_01v8 ad=1.25e+11p pd=1.5e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=7.2e+11p pd=5.44e+06u as=3.9e+11p ps=2.78e+06u w=1e+06u l=150000u
X2 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B a_94_6# GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=0p ps=0u w=500000u l=150000u
.ends

.subckt inv VDD GND Y A
X0 Y A GND GND sky130_fd_pr__nfet_01v8 ad=1.8e+11p pd=1.72e+06u as=1.8e+11p ps=1.72e+06u w=500000u l=150000u
X1 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=3.6e+11p pd=2.72e+06u as=3.6e+11p ps=2.72e+06u w=1e+06u l=150000u
.ends

*.subckt multiplexor A2 Y2 B2 A3 Y3 B3 A0 Y0 B0 A1 Y1 B1 A6 Y6 B6 A7 Y7 B7 A4 Y4 B4
+ A5 Y5 B5 SEL
Xnand2_18 VDD GND nand2_19/A A6 SEL nand2
Xnand2_6 VDD GND nand2_7/A A2 SEL nand2
Xnand2_19 VDD GND Y6 nand2_19/A nand2_21/Y nand2
Xnand2_7 VDD GND Y2 nand2_7/A nand2_8/Y nand2
Xnand2_8 VDD GND nand2_8/Y inv_0/Y B2 nand2
Xnand2_9 VDD GND nand2_9/Y A3 SEL nand2
Xinv_0 VDD GND inv_0/Y SEL inv
Xnand2_20 VDD GND nand2_22/A A7 SEL nand2
Xnand2_21 VDD GND nand2_21/Y inv_0/Y B6 nand2
Xnand2_10 VDD GND Y3 nand2_9/Y nand2_11/Y nand2
Xnand2_22 VDD GND Y7 nand2_22/A nand2_23/Y nand2
Xnand2_11 VDD GND nand2_11/Y inv_0/Y B3 nand2
Xnand2_23 VDD GND nand2_23/Y inv_0/Y B7 nand2
Xnand2_12 VDD GND nand2_13/A A4 SEL nand2
Xnand2_0 VDD GND nand2_1/A A0 SEL nand2
Xnand2_13 VDD GND Y4 nand2_13/A nand2_14/Y nand2
Xnand2_2 VDD GND nand2_2/Y inv_0/Y B0 nand2
Xnand2_1 VDD GND Y0 nand2_1/A nand2_2/Y nand2
Xnand2_14 VDD GND nand2_14/Y inv_0/Y B4 nand2
Xnand2_3 VDD GND nand2_4/B inv_0/Y B1 nand2
Xnand2_16 VDD GND Y5 nand2_16/A nand2_17/Y nand2
Xnand2_15 VDD GND nand2_16/A A5 SEL nand2
Xnand2_4 VDD GND Y1 nand2_5/Y nand2_4/B nand2
Xnand2_17 VDD GND nand2_17/Y inv_0/Y B5 nand2
Xnand2_5 VDD GND nand2_5/Y A1 SEL nand2
*.ends

