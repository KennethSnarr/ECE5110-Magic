magic
tech sky130A
timestamp 1677803710
<< nwell >>
rect -42 135 157 426
<< nmos >>
rect 32 3 47 53
rect 68 3 83 53
<< pmos >>
rect 32 253 47 353
rect 68 253 83 353
<< ndiff >>
rect -4 45 32 53
rect -4 11 4 45
rect 21 11 32 45
rect -4 3 32 11
rect 47 3 68 53
rect 83 45 119 53
rect 83 11 94 45
rect 111 11 119 45
rect 83 3 119 11
<< pdiff >>
rect -4 345 32 353
rect -4 261 4 345
rect 21 261 32 345
rect -4 253 32 261
rect 47 253 68 353
rect 83 345 119 353
rect 83 261 94 345
rect 111 261 119 345
rect 83 253 119 261
<< ndiffc >>
rect 4 11 21 45
rect 94 11 111 45
<< pdiffc >>
rect 4 261 21 345
rect 94 261 111 345
<< psubdiff >>
rect -4 -52 8 -24
rect 111 -52 123 -24
<< nsubdiff >>
rect 3 380 15 408
rect 118 380 130 408
<< psubdiffcont >>
rect 8 -52 111 -24
<< nsubdiffcont >>
rect 15 380 118 408
<< poly >>
rect 32 353 47 366
rect 68 353 83 366
rect 32 170 47 253
rect 68 209 83 253
rect 68 201 149 209
rect 68 194 124 201
rect 116 184 124 194
rect 141 184 149 201
rect 116 176 149 184
rect -1 162 47 170
rect -1 145 7 162
rect 24 145 47 162
rect -1 137 47 145
rect 32 53 47 137
rect 116 125 149 133
rect 116 115 124 125
rect 68 108 124 115
rect 141 108 149 125
rect 68 100 149 108
rect 68 53 83 100
rect 32 -10 47 3
rect 68 -10 83 3
<< polycont >>
rect 124 184 141 201
rect 7 145 24 162
rect 124 108 141 125
<< locali >>
rect -40 408 155 418
rect -40 380 15 408
rect 118 380 155 408
rect -40 370 155 380
rect -4 345 29 370
rect -4 261 4 345
rect 21 261 29 345
rect -4 253 29 261
rect 86 345 119 353
rect 86 261 94 345
rect 111 261 119 345
rect 86 243 119 261
rect 50 226 119 243
rect -1 162 32 170
rect -1 145 7 162
rect 24 145 32 162
rect -1 137 32 145
rect 50 81 68 226
rect 116 201 149 209
rect 116 184 124 201
rect 141 184 149 201
rect 116 176 149 184
rect 116 125 149 133
rect 116 108 124 125
rect 141 108 149 125
rect 116 100 149 108
rect 50 64 119 81
rect -4 45 29 53
rect -4 11 4 45
rect 21 11 29 45
rect -4 -14 29 11
rect 86 45 119 64
rect 86 11 94 45
rect 111 11 119 45
rect 86 3 119 11
rect -40 -24 155 -14
rect -40 -52 8 -24
rect 111 -52 155 -24
rect -40 -62 155 -52
<< labels >>
flabel locali -1 137 32 170 0 FreeSerif 80 0 0 0 A
port 7 nsew
flabel nwell -40 370 156 418 0 FreeSerif 80 0 0 0 VDD!
port 0 nsew
flabel locali 116 100 149 133 0 FreeSerif 80 0 0 0 EN
port 8 nsew
flabel locali 116 176 149 209 0 FreeSerif 80 0 0 0 NOT_EN
port 9 nsew
flabel locali -40 -62 155 -14 0 FreeSerif 80 0 0 0 GND!
port 1 nsew
<< end >>
