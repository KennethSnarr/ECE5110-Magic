magic
tech sky130A
timestamp 1679435600
<< nwell >>
rect -42 135 793 426
<< nmos >>
rect 32 3 47 53
rect 72 3 87 53
rect 200 3 215 53
rect 240 3 255 53
rect 368 3 383 53
rect 482 3 497 53
rect 522 3 537 53
rect 650 3 665 53
rect 690 3 705 53
<< pmos >>
rect 32 253 47 353
rect 86 253 101 353
rect 200 253 215 353
rect 254 253 269 353
rect 368 253 383 353
rect 482 253 497 353
rect 536 253 551 353
rect 650 253 665 353
rect 704 253 719 353
<< ndiff >>
rect -4 45 32 53
rect -4 11 4 45
rect 21 11 32 45
rect -4 3 32 11
rect 47 3 72 53
rect 87 45 123 53
rect 87 11 98 45
rect 115 11 123 45
rect 87 3 123 11
rect 164 45 200 53
rect 164 11 172 45
rect 189 11 200 45
rect 164 3 200 11
rect 215 3 240 53
rect 255 45 291 53
rect 255 11 266 45
rect 283 11 291 45
rect 255 3 291 11
rect 332 45 368 53
rect 332 11 340 45
rect 357 11 368 45
rect 332 3 368 11
rect 383 45 419 53
rect 383 11 394 45
rect 411 11 419 45
rect 383 3 419 11
rect 446 45 482 53
rect 446 11 454 45
rect 471 11 482 45
rect 446 3 482 11
rect 497 3 522 53
rect 537 45 573 53
rect 537 11 548 45
rect 565 11 573 45
rect 537 3 573 11
rect 614 45 650 53
rect 614 11 622 45
rect 639 11 650 45
rect 614 3 650 11
rect 665 3 690 53
rect 705 45 741 53
rect 705 11 716 45
rect 733 11 741 45
rect 705 3 741 11
<< pdiff >>
rect -4 345 32 353
rect -4 261 4 345
rect 21 261 32 345
rect -4 253 32 261
rect 47 345 86 353
rect 47 261 58 345
rect 75 261 86 345
rect 47 253 86 261
rect 101 345 137 353
rect 101 261 112 345
rect 129 261 137 345
rect 101 253 137 261
rect 164 345 200 353
rect 164 261 172 345
rect 189 261 200 345
rect 164 253 200 261
rect 215 345 254 353
rect 215 261 226 345
rect 243 261 254 345
rect 215 253 254 261
rect 269 345 305 353
rect 269 261 280 345
rect 297 261 305 345
rect 269 253 305 261
rect 332 345 368 353
rect 332 261 340 345
rect 357 261 368 345
rect 332 253 368 261
rect 383 345 419 353
rect 383 261 394 345
rect 411 261 419 345
rect 383 253 419 261
rect 446 345 482 353
rect 446 261 454 345
rect 471 261 482 345
rect 446 253 482 261
rect 497 345 536 353
rect 497 261 508 345
rect 525 261 536 345
rect 497 253 536 261
rect 551 345 587 353
rect 551 261 562 345
rect 579 261 587 345
rect 551 253 587 261
rect 614 345 650 353
rect 614 261 622 345
rect 639 261 650 345
rect 614 253 650 261
rect 665 345 704 353
rect 665 261 676 345
rect 693 261 704 345
rect 665 253 704 261
rect 719 345 755 353
rect 719 261 730 345
rect 747 261 755 345
rect 719 253 755 261
<< ndiffc >>
rect 4 11 21 45
rect 98 11 115 45
rect 172 11 189 45
rect 266 11 283 45
rect 340 11 357 45
rect 394 11 411 45
rect 454 11 471 45
rect 548 11 565 45
rect 622 11 639 45
rect 716 11 733 45
<< pdiffc >>
rect 4 261 21 345
rect 58 261 75 345
rect 112 261 129 345
rect 172 261 189 345
rect 226 261 243 345
rect 280 261 297 345
rect 340 261 357 345
rect 394 261 411 345
rect 454 261 471 345
rect 508 261 525 345
rect 562 261 579 345
rect 622 261 639 345
rect 676 261 693 345
rect 730 261 747 345
<< psubdiff >>
rect -4 -52 8 -24
rect 729 -52 741 -24
<< nsubdiff >>
rect -4 380 8 408
rect 743 380 755 408
<< psubdiffcont >>
rect 8 -52 729 -24
<< nsubdiffcont >>
rect 8 380 743 408
<< poly >>
rect 32 353 47 366
rect 86 353 101 366
rect 200 353 215 366
rect 254 353 269 366
rect 368 353 383 366
rect 482 353 497 366
rect 536 353 551 366
rect 650 353 665 366
rect 704 353 719 366
rect 32 235 47 253
rect -1 227 47 235
rect -1 210 7 227
rect 24 210 47 227
rect -1 202 47 210
rect 32 53 47 202
rect 86 185 101 253
rect 200 185 215 253
rect 86 177 215 185
rect 86 160 141 177
rect 158 160 215 177
rect 86 152 215 160
rect 86 99 101 152
rect 72 84 101 99
rect 72 53 87 84
rect 200 53 215 152
rect 254 185 269 253
rect 368 235 383 253
rect 335 227 383 235
rect 335 210 343 227
rect 360 210 383 227
rect 335 202 383 210
rect 254 177 302 185
rect 254 160 277 177
rect 294 160 302 177
rect 254 152 302 160
rect 254 99 269 152
rect 240 84 269 99
rect 240 53 255 84
rect 368 53 383 202
rect 482 170 497 253
rect 449 162 497 170
rect 449 145 457 162
rect 474 145 497 162
rect 449 137 497 145
rect 482 53 497 137
rect 536 211 551 253
rect 536 203 584 211
rect 536 186 559 203
rect 576 186 584 203
rect 536 178 584 186
rect 536 99 551 178
rect 650 170 665 253
rect 617 162 665 170
rect 617 145 625 162
rect 642 145 665 162
rect 617 137 665 145
rect 522 84 551 99
rect 522 53 537 84
rect 650 53 665 137
rect 704 211 719 253
rect 704 203 752 211
rect 704 186 727 203
rect 744 186 752 203
rect 704 178 752 186
rect 704 99 719 178
rect 690 84 719 99
rect 690 53 705 84
rect 32 -10 47 3
rect 72 -10 87 3
rect 200 -10 215 3
rect 240 -10 255 3
rect 368 -10 383 3
rect 482 -10 497 3
rect 522 -10 537 3
rect 650 -10 665 3
rect 690 -10 705 3
<< polycont >>
rect 7 210 24 227
rect 141 160 158 177
rect 343 210 360 227
rect 277 160 294 177
rect 457 145 474 162
rect 559 186 576 203
rect 625 145 642 162
rect 727 186 744 203
<< locali >>
rect -40 408 791 418
rect -40 380 8 408
rect 743 380 791 408
rect -40 370 791 380
rect -4 345 29 370
rect -4 261 4 345
rect 21 261 29 345
rect -4 253 29 261
rect 50 345 83 353
rect 50 261 58 345
rect 75 261 83 345
rect -1 227 32 235
rect -1 210 7 227
rect 24 210 32 227
rect -1 202 32 210
rect 50 135 83 261
rect 104 345 137 370
rect 104 261 112 345
rect 129 261 137 345
rect 104 253 137 261
rect 164 345 197 370
rect 164 261 172 345
rect 189 261 197 345
rect 164 253 197 261
rect 218 345 251 353
rect 218 261 226 345
rect 243 261 251 345
rect 101 177 200 185
rect 101 160 141 177
rect 158 160 200 177
rect 101 152 200 160
rect 218 135 251 261
rect 272 345 305 370
rect 272 261 280 345
rect 297 261 305 345
rect 272 253 305 261
rect 332 345 365 370
rect 332 261 340 345
rect 357 261 365 345
rect 332 253 365 261
rect 386 345 419 353
rect 386 261 394 345
rect 411 261 419 345
rect 335 227 368 235
rect 335 210 343 227
rect 360 210 368 227
rect 335 202 368 210
rect 269 177 302 185
rect 269 160 277 177
rect 294 160 302 177
rect 269 152 302 160
rect 386 177 419 261
rect 446 345 479 370
rect 446 261 454 345
rect 471 261 479 345
rect 446 253 479 261
rect 500 345 533 353
rect 500 261 508 345
rect 525 261 533 345
rect 386 160 394 177
rect 411 160 419 177
rect 50 127 156 135
rect 50 110 131 127
rect 148 110 156 127
rect 50 102 156 110
rect 218 102 291 135
rect -4 45 29 53
rect -4 11 4 45
rect 21 11 29 45
rect -4 -14 29 11
rect 90 45 123 102
rect 258 77 291 102
rect 258 60 266 77
rect 283 60 291 77
rect 90 11 98 45
rect 115 11 123 45
rect 90 3 123 11
rect 164 45 197 53
rect 164 11 172 45
rect 189 11 197 45
rect 164 -14 197 11
rect 258 45 291 60
rect 258 11 266 45
rect 283 11 291 45
rect 258 3 291 11
rect 332 45 365 53
rect 332 11 340 45
rect 357 11 365 45
rect 332 -14 365 11
rect 386 45 419 160
rect 449 162 482 170
rect 449 145 457 162
rect 474 145 482 162
rect 449 137 482 145
rect 500 162 533 261
rect 554 345 587 370
rect 554 261 562 345
rect 579 261 587 345
rect 554 253 587 261
rect 614 345 647 370
rect 614 261 622 345
rect 639 261 647 345
rect 614 253 647 261
rect 668 345 701 353
rect 668 261 676 345
rect 693 261 701 345
rect 551 203 584 211
rect 551 186 559 203
rect 576 186 584 203
rect 551 178 584 186
rect 668 203 701 261
rect 722 345 755 370
rect 722 261 730 345
rect 747 261 755 345
rect 722 253 755 261
rect 668 186 676 203
rect 693 186 701 203
rect 500 145 508 162
rect 525 145 533 162
rect 500 135 533 145
rect 617 162 650 170
rect 617 145 625 162
rect 642 145 650 162
rect 617 137 650 145
rect 668 135 701 186
rect 719 203 752 211
rect 719 186 727 203
rect 744 186 752 203
rect 719 178 752 186
rect 500 102 573 135
rect 668 102 741 135
rect 386 11 394 45
rect 411 11 419 45
rect 386 3 419 11
rect 446 45 479 53
rect 446 11 454 45
rect 471 11 479 45
rect 446 -14 479 11
rect 540 45 573 102
rect 540 11 548 45
rect 565 11 573 45
rect 540 3 573 11
rect 614 45 647 53
rect 614 11 622 45
rect 639 11 647 45
rect 614 -14 647 11
rect 708 45 741 102
rect 708 11 716 45
rect 733 11 741 45
rect 708 3 741 11
rect -40 -24 791 -14
rect -40 -52 8 -24
rect 729 -52 791 -24
rect -40 -62 791 -52
<< viali >>
rect 7 210 24 227
rect 343 210 360 227
rect 277 160 294 177
rect 394 160 411 177
rect 131 110 148 127
rect 266 60 283 77
rect 457 145 474 162
rect 559 186 576 203
rect 676 186 693 203
rect 508 145 525 162
rect 625 145 642 162
rect 727 186 744 203
<< metal1 >>
rect -1 227 368 235
rect -1 210 7 227
rect 24 220 343 227
rect 24 210 32 220
rect -1 202 32 210
rect 335 210 343 220
rect 360 210 368 227
rect 335 202 368 210
rect 551 203 584 211
rect 668 203 701 211
rect 551 186 559 203
rect 576 186 676 203
rect 693 186 701 203
rect 269 177 302 185
rect 386 177 419 185
rect 551 178 584 186
rect 668 178 701 186
rect 719 203 752 211
rect 719 186 727 203
rect 744 186 752 203
rect 719 178 752 186
rect 269 160 277 177
rect 294 160 394 177
rect 411 160 419 177
rect 269 152 302 160
rect 386 152 419 160
rect 449 162 482 170
rect 449 145 457 162
rect 474 145 482 162
rect 449 137 482 145
rect 500 162 533 170
rect 617 162 650 170
rect 500 145 508 162
rect 525 145 625 162
rect 642 145 650 162
rect 500 137 533 145
rect 617 137 650 145
rect 123 127 156 135
rect 123 110 131 127
rect 148 126 156 127
rect 449 126 474 137
rect 148 110 474 126
rect 727 122 744 178
rect 123 102 156 110
rect 490 107 744 122
rect 258 77 291 83
rect 490 77 504 107
rect 258 60 266 77
rect 283 62 504 77
rect 283 60 291 62
rect 258 53 291 60
<< labels >>
flabel locali -40 -62 791 -14 0 FreeSerif 80 0 0 0 GND!
port 11 nsew
flabel locali -40 370 791 418 0 FreeSerif 80 0 0 0 VDD!
port 0 nsew
flabel locali s -1 202 32 235 0 FreeSerif 80 0 0 0 D
port 1 nsew
flabel locali s 101 152 200 185 0 FreeSerif 80 0 0 0 CLK
port 6 nsew
flabel locali s 540 53 573 135 0 FreeSerif 80 0 0 0 Q
port 22 nsew
flabel locali s 708 53 741 135 0 FreeSerif 80 0 0 0 NOT_Q
port 23 nsew
rlabel ndiff 32 24 32 24 0 S$
rlabel ndiff 72 24 72 24 0 S$
rlabel ndiff 200 24 200 24 0 S$
rlabel ndiff 240 24 240 24 0 S$
rlabel ndiff 368 24 368 24 0 S$
rlabel ndiff 482 22 482 22 0 S$
rlabel ndiff 522 22 522 22 0 S$
rlabel ndiff 650 20 650 20 0 S$
rlabel ndiff 690 18 690 18 0 S$
rlabel pdiff 719 312 719 312 0 S$
rlabel pdiff 650 310 650 310 0 S$
rlabel pdiff 551 314 551 314 0 S$
rlabel pdiff 482 312 482 312 0 S$
rlabel pdiff 368 318 368 318 0 S$
rlabel pdiff 269 314 269 314 0 S$
rlabel pdiff 200 320 200 320 0 S$
rlabel pdiff 101 312 101 312 0 S$
rlabel pdiff 32 314 32 314 0 S$
<< end >>
