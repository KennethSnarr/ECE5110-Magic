magic
tech sky130A
magscale 1 2
timestamp 1682034221
<< locali >>
rect -222 910 18748 1006
rect -222 -722 -126 910
rect 367 574 382 640
rect 3768 574 3781 640
rect 316 572 382 574
rect 48 442 114 510
rect 10404 444 10470 510
rect 10672 498 10738 510
rect 10672 458 10694 498
rect 10734 458 10738 498
rect 10672 444 10738 458
rect 2970 325 3036 440
rect 2970 276 3036 283
rect 3306 311 3372 440
rect 3306 276 3372 277
rect 6422 326 6488 440
rect 6422 276 6488 277
rect 6758 314 6824 440
rect 9874 308 9940 440
rect 10210 326 10276 440
rect 11110 374 11176 676
rect 11548 571 11614 592
rect 11680 499 11746 510
rect 11680 459 11686 499
rect 11726 459 11746 499
rect 11680 444 11746 459
rect 12118 374 12184 676
rect 12556 584 12622 592
rect 12556 544 12578 584
rect 12618 544 12622 584
rect 12556 526 12622 544
rect 12688 501 12754 510
rect 12688 461 12696 501
rect 12736 461 12754 501
rect 12688 444 12754 461
rect 13126 374 13192 676
rect 13564 567 13630 592
rect 13696 501 13762 510
rect 13696 461 13700 501
rect 13740 461 13762 501
rect 13696 444 13762 461
rect 14134 374 14200 676
rect 14572 580 14638 592
rect 14572 540 14576 580
rect 14616 540 14638 580
rect 14572 526 14638 540
rect 14704 497 14770 510
rect 14704 457 14714 497
rect 14754 457 14770 497
rect 14704 444 14770 457
rect 15142 374 15208 676
rect 15580 564 15646 592
rect 15712 499 15778 510
rect 15712 459 15720 499
rect 15760 459 15778 499
rect 15712 444 15778 459
rect 16150 374 16216 676
rect 16588 580 16654 592
rect 16588 540 16600 580
rect 16640 540 16654 580
rect 16588 526 16654 540
rect 16720 503 16786 510
rect 16720 463 16726 503
rect 16766 463 16786 503
rect 16720 444 16786 463
rect 17158 374 17224 676
rect 17596 566 17662 592
rect 17728 497 17794 510
rect 17728 457 17736 497
rect 17776 457 17794 497
rect 17728 444 17794 457
rect 18166 374 18232 676
rect 18604 573 18670 592
rect 18604 539 18609 573
rect 18643 539 18670 573
rect 18604 526 18670 539
rect 10210 263 10276 276
rect -30 46 18748 142
rect 2970 -89 3036 -88
rect 2970 -252 3036 -130
rect 3306 -252 3372 -138
rect 6422 -252 6488 -134
rect 6758 -252 6824 -133
rect 48 -322 114 -256
rect 3500 -322 3566 -256
rect 316 -452 382 -386
rect 3768 -452 3834 -386
rect -222 -818 15296 -722
rect -222 -2450 -126 -818
rect 316 -1154 332 -1088
rect 3768 -1156 3834 -1140
rect 6952 -1284 7018 -1218
rect 7220 -1236 7286 -1218
rect 7220 -1276 7233 -1236
rect 7273 -1276 7286 -1236
rect 7220 -1284 7286 -1276
rect 7658 -1288 7724 -1052
rect 8096 -1202 8162 -1177
rect 8228 -1234 8294 -1218
rect 8228 -1274 8235 -1234
rect 8275 -1274 8294 -1234
rect 8228 -1284 8294 -1274
rect 8666 -1265 8732 -1052
rect 9104 -1161 9170 -1136
rect 2970 -1404 3036 -1288
rect 3306 -1400 3372 -1288
rect 3306 -1452 3372 -1451
rect 6422 -1416 6488 -1288
rect 6758 -1406 6824 -1288
rect 7658 -1354 7724 -1336
rect 9236 -1232 9302 -1218
rect 9236 -1272 9247 -1232
rect 9287 -1272 9302 -1232
rect 9236 -1284 9302 -1272
rect 9674 -1253 9740 -1052
rect 10112 -1159 10178 -1136
rect 8666 -1354 8732 -1306
rect 9674 -1293 9692 -1253
rect 9732 -1293 9740 -1253
rect 10244 -1234 10310 -1218
rect 10244 -1274 10260 -1234
rect 10300 -1274 10310 -1234
rect 10244 -1284 10310 -1274
rect 10682 -1257 10748 -1052
rect 11120 -1150 11186 -1136
rect 11120 -1162 11132 -1150
rect 11180 -1162 11186 -1150
rect 9674 -1354 9740 -1293
rect 11252 -1230 11318 -1218
rect 11252 -1270 11266 -1230
rect 11306 -1270 11318 -1230
rect 11252 -1284 11318 -1270
rect 11690 -1254 11756 -1052
rect 12128 -1143 12194 -1136
rect 12128 -1183 12145 -1143
rect 12185 -1183 12194 -1143
rect 12128 -1202 12194 -1183
rect 10682 -1354 10748 -1295
rect 11690 -1294 11700 -1254
rect 11734 -1294 11756 -1254
rect 12260 -1232 12326 -1218
rect 12260 -1272 12281 -1232
rect 12321 -1272 12326 -1232
rect 12260 -1284 12326 -1272
rect 12698 -1269 12764 -1052
rect 13136 -1152 13202 -1136
rect 13136 -1192 13148 -1152
rect 13188 -1192 13202 -1152
rect 13136 -1202 13202 -1192
rect 11690 -1354 11756 -1294
rect 13268 -1228 13334 -1218
rect 13268 -1268 13280 -1228
rect 13320 -1268 13334 -1228
rect 13268 -1284 13334 -1268
rect 13706 -1242 13772 -1052
rect 14714 -1083 14780 -1052
rect 14144 -1143 14210 -1136
rect 14144 -1183 14148 -1143
rect 14188 -1183 14210 -1143
rect 14144 -1202 14210 -1183
rect 13706 -1282 13714 -1242
rect 13754 -1282 13772 -1242
rect 12698 -1354 12764 -1307
rect 13706 -1354 13772 -1282
rect 14276 -1234 14342 -1218
rect 14276 -1274 14295 -1234
rect 14335 -1274 14342 -1234
rect 14276 -1284 14342 -1274
rect 14714 -1354 14780 -1123
rect 15152 -1142 15218 -1136
rect 15152 -1182 15178 -1142
rect 15152 -1202 15218 -1182
rect 15546 -1586 15642 46
rect -30 -1682 15642 -1586
rect 2970 -1980 3036 -1877
rect 3306 -1817 3372 -1816
rect 3306 -1980 3372 -1864
rect 6422 -1980 6488 -1864
rect 6758 -1821 6824 -1816
rect 6758 -1980 6824 -1872
rect 6952 -2050 7018 -1933
rect 7658 -1979 7724 -1914
rect 7220 -2050 7286 -2034
rect 8666 -1979 8732 -1914
rect 3768 -2180 3774 -2114
rect 7658 -2216 7724 -2028
rect 8228 -2001 8294 -1984
rect 8228 -2041 8238 -2001
rect 8278 -2041 8294 -2001
rect 8228 -2050 8294 -2041
rect 9674 -1945 9740 -1914
rect 8096 -2082 8162 -2066
rect 8096 -2122 8120 -2082
rect 8160 -2122 8162 -2082
rect 8096 -2132 8162 -2122
rect 8666 -2216 8732 -2041
rect 9236 -1998 9302 -1984
rect 9236 -2038 9246 -1998
rect 9286 -2038 9302 -1998
rect 9236 -2050 9302 -2038
rect 10682 -1969 10748 -1914
rect 9104 -2082 9170 -2066
rect 9104 -2122 9110 -2082
rect 9150 -2122 9170 -2082
rect 9104 -2132 9170 -2122
rect 9674 -2216 9740 -1986
rect 10244 -1995 10310 -1984
rect 10244 -2035 10252 -1995
rect 10292 -2035 10310 -1995
rect 10244 -2050 10310 -2035
rect 11690 -1963 11756 -1914
rect 10112 -2078 10178 -2066
rect 10112 -2118 10120 -2078
rect 10160 -2118 10178 -2078
rect 10112 -2132 10178 -2118
rect 10682 -2216 10748 -2013
rect 11252 -2002 11318 -1984
rect 11252 -2042 11258 -2002
rect 11298 -2042 11318 -2002
rect 11252 -2050 11318 -2042
rect 12698 -1963 12764 -1914
rect 11120 -2079 11186 -2066
rect 11120 -2119 11138 -2079
rect 11178 -2119 11186 -2079
rect 11120 -2132 11186 -2119
rect 11690 -2216 11756 -2007
rect 12260 -1993 12326 -1984
rect 12260 -2033 12268 -1993
rect 12308 -2033 12326 -1993
rect 12260 -2050 12326 -2033
rect 13706 -1967 13772 -1914
rect 12128 -2080 12194 -2066
rect 12128 -2120 12146 -2080
rect 12186 -2120 12194 -2080
rect 12128 -2132 12194 -2120
rect 12698 -2216 12764 -2000
rect 13268 -2000 13334 -1984
rect 13268 -2040 13274 -2000
rect 13314 -2040 13334 -2000
rect 13268 -2050 13334 -2040
rect 14714 -1973 14780 -1914
rect 13136 -2088 13202 -2066
rect 13136 -2128 13150 -2088
rect 13190 -2128 13202 -2088
rect 13136 -2132 13202 -2128
rect 13706 -2216 13772 -2007
rect 14276 -1993 14342 -1984
rect 14276 -2033 14286 -1993
rect 14326 -2033 14342 -1993
rect 14276 -2050 14342 -2033
rect 14144 -2075 14210 -2066
rect 14144 -2115 14157 -2075
rect 14197 -2115 14210 -2075
rect 14144 -2132 14210 -2115
rect 14714 -2216 14780 -2018
rect 15152 -2132 15218 -2106
rect -222 -2546 15296 -2450
<< viali >>
rect 316 574 367 640
rect 3781 574 3834 640
rect 7220 574 7286 640
rect 3500 444 3566 510
rect 6952 444 7018 510
rect 10694 458 10734 498
rect 2970 283 3036 325
rect 3306 277 3372 311
rect 6422 277 6488 326
rect 6758 265 6824 314
rect 9874 265 9940 308
rect 11548 526 11614 571
rect 11686 459 11726 499
rect 12578 544 12618 584
rect 12696 461 12736 501
rect 13564 526 13630 567
rect 13700 461 13740 501
rect 14576 540 14616 580
rect 14714 457 14754 497
rect 15580 526 15646 564
rect 15720 459 15760 499
rect 16600 540 16640 580
rect 16726 463 16766 503
rect 17596 526 17662 566
rect 17736 457 17776 497
rect 18609 539 18643 573
rect 10210 276 10276 326
rect 2970 -130 3036 -89
rect 3306 -138 3372 -87
rect 6422 -134 6488 -85
rect 6758 -133 6824 -83
rect 332 -1154 382 -1088
rect 3768 -1140 3834 -1088
rect 48 -1284 114 -1218
rect 3500 -1284 3566 -1218
rect 7233 -1276 7273 -1236
rect 8096 -1177 8162 -1136
rect 8235 -1274 8275 -1234
rect 9104 -1202 9170 -1161
rect 2970 -1457 3036 -1404
rect 3306 -1451 3372 -1400
rect 6422 -1467 6488 -1416
rect 7658 -1336 7724 -1288
rect 8666 -1306 8732 -1265
rect 9247 -1272 9287 -1232
rect 10112 -1202 10178 -1159
rect 9692 -1293 9732 -1253
rect 10260 -1274 10300 -1234
rect 11132 -1162 11180 -1150
rect 11120 -1202 11186 -1162
rect 10682 -1295 10748 -1257
rect 11266 -1270 11306 -1230
rect 12145 -1183 12185 -1143
rect 11700 -1294 11734 -1254
rect 12281 -1272 12321 -1232
rect 13148 -1192 13188 -1152
rect 12698 -1307 12764 -1269
rect 13280 -1268 13320 -1228
rect 14714 -1123 14780 -1083
rect 14148 -1183 14188 -1143
rect 13714 -1282 13754 -1242
rect 14295 -1274 14335 -1234
rect 15178 -1182 15218 -1142
rect 6758 -1459 6824 -1406
rect 2970 -1877 3036 -1811
rect 3306 -1864 3372 -1817
rect 6422 -1864 6488 -1815
rect 6758 -1872 6824 -1821
rect 6952 -1933 7018 -1899
rect 48 -2050 114 -1984
rect 3500 -2050 3566 -1984
rect 7220 -2034 7286 -1984
rect 7658 -2028 7724 -1979
rect 316 -2180 382 -2114
rect 3774 -2180 3834 -2114
rect 8238 -2041 8278 -2001
rect 8666 -2041 8732 -1979
rect 8120 -2122 8160 -2082
rect 9246 -2038 9286 -1998
rect 9674 -1986 9740 -1945
rect 9110 -2122 9150 -2082
rect 10252 -2035 10292 -1995
rect 10682 -2013 10748 -1969
rect 10120 -2118 10160 -2078
rect 11258 -2042 11298 -2002
rect 11690 -2007 11756 -1963
rect 11138 -2119 11178 -2079
rect 12268 -2033 12308 -1993
rect 12698 -2000 12764 -1963
rect 12146 -2120 12186 -2080
rect 13274 -2040 13314 -2000
rect 13706 -2007 13772 -1967
rect 13150 -2128 13190 -2088
rect 14286 -2033 14326 -1993
rect 14714 -2018 14780 -1973
rect 14157 -2115 14197 -2075
rect 15152 -2106 15218 -2066
<< metal1 >>
rect 10211 991 10217 992
rect 7223 941 10217 991
rect 310 640 373 652
rect 310 632 316 640
rect 302 580 308 632
rect 310 574 316 580
rect 367 574 373 640
rect 310 562 373 574
rect 3775 640 3840 652
rect 7223 646 7273 941
rect 10211 940 10217 941
rect 10269 940 10275 992
rect 3775 574 3781 640
rect 3834 574 3840 640
rect 3775 562 3840 574
rect 7208 640 7298 646
rect 7208 574 7220 640
rect 7286 574 7298 640
rect 11542 577 11620 578
rect 7208 568 7298 574
rect 11536 572 11626 577
rect 3494 510 3572 522
rect 11536 520 11542 572
rect 11620 520 11626 572
rect 12566 538 12572 590
rect 12624 538 12630 590
rect 13558 573 13636 578
rect 13552 572 13642 573
rect 13552 520 13558 572
rect 13636 520 13642 572
rect 14564 534 14570 586
rect 14622 534 14628 586
rect 15574 571 15652 577
rect 15568 520 15574 570
rect 3494 444 3500 510
rect 3566 444 3572 510
rect 3494 432 3572 444
rect 6940 510 7030 516
rect 11542 514 11620 520
rect 13558 514 13636 520
rect 15652 520 15658 570
rect 16588 534 16594 586
rect 16646 534 16652 586
rect 17590 572 17668 578
rect 18603 573 18649 585
rect 17584 520 17590 572
rect 17668 520 17674 572
rect 18603 539 18609 573
rect 18643 539 18649 573
rect 18603 527 18649 539
rect 15574 513 15652 519
rect 17590 514 17668 520
rect 6940 444 6952 510
rect 7018 494 7030 510
rect 6940 442 6970 444
rect 7022 442 7030 494
rect 10682 452 10688 504
rect 10740 452 10746 504
rect 11674 453 11680 505
rect 11732 453 11738 505
rect 12684 455 12690 507
rect 12742 455 12748 507
rect 13688 455 13694 507
rect 13746 455 13752 507
rect 14702 451 14708 503
rect 14760 451 14766 503
rect 15708 453 15714 505
rect 15766 453 15772 505
rect 16714 457 16720 509
rect 16772 457 16778 509
rect 17724 451 17730 503
rect 17782 451 17788 503
rect 6940 438 7030 442
rect 6970 436 7022 438
rect -41 329 -35 381
rect 17 329 23 381
rect -27 -2512 8 329
rect 2958 325 3048 331
rect 2958 283 2970 325
rect 3036 283 3048 325
rect 3300 320 3378 326
rect 2958 277 3048 283
rect 2982 186 3024 277
rect 3294 271 3300 317
rect 3378 271 3384 317
rect 3300 262 3378 268
rect 2977 180 3029 186
rect 2977 125 3029 128
rect 54 122 3029 125
rect 54 111 3024 122
rect 3504 120 3553 432
rect 10204 332 10282 338
rect 6410 326 6500 332
rect 6410 323 6422 326
rect 6488 323 6500 326
rect 6410 271 6416 323
rect 6494 271 6500 323
rect 6746 314 6836 320
rect 9868 314 9946 317
rect 6746 311 6758 314
rect 6824 311 6836 314
rect 6416 265 6494 271
rect 6746 259 6752 311
rect 6830 259 6836 311
rect 9862 311 9952 314
rect 9862 259 9868 311
rect 9946 259 9952 311
rect 10198 280 10204 332
rect 10282 280 10288 332
rect 10198 276 10210 280
rect 10276 276 10288 280
rect 10198 270 10288 276
rect 6752 253 6830 259
rect 9868 253 9946 259
rect 54 88 3022 111
rect 54 -320 91 88
rect 3504 71 6480 120
rect 6431 11 6480 71
rect 11906 25 11958 31
rect 15006 28 15066 34
rect 11546 20 11552 22
rect 6431 -39 7002 11
rect 2964 -83 3042 -77
rect 3300 -81 3378 -75
rect 6431 -79 6480 -39
rect 2958 -135 2964 -83
rect 3042 -135 3048 -83
rect 2958 -136 3048 -135
rect 3294 -133 3300 -81
rect 3378 -133 3384 -81
rect 2964 -141 3042 -136
rect 3294 -138 3306 -133
rect 3372 -138 3384 -133
rect 3294 -144 3384 -138
rect 6410 -85 6500 -79
rect 6410 -134 6422 -85
rect 6488 -134 6500 -85
rect 6410 -140 6500 -134
rect 6746 -83 6836 -77
rect 6746 -87 6758 -83
rect 6824 -87 6836 -83
rect 6746 -139 6752 -87
rect 6830 -139 6836 -87
rect 6952 -138 7002 -39
rect 7667 -28 11552 20
rect 6752 -145 6830 -139
rect 6945 -190 6951 -138
rect 7003 -190 7009 -138
rect 321 -445 327 -393
rect 379 -445 385 -393
rect 3511 -747 3562 -257
rect 3776 -440 3782 -388
rect 3834 -440 3840 -388
rect 6650 -604 6702 -598
rect 3670 -658 3676 -606
rect 3728 -611 3734 -606
rect 3884 -611 3890 -605
rect 3728 -652 3890 -611
rect 3728 -658 3734 -652
rect 3884 -657 3890 -652
rect 3942 -657 3948 -605
rect 6702 -650 6916 -609
rect 6650 -662 6702 -656
rect 6875 -737 6916 -650
rect 3511 -798 6482 -747
rect 6864 -789 6870 -737
rect 6922 -789 6928 -737
rect 6431 -912 6482 -798
rect 7667 -884 7715 -28
rect 11546 -30 11552 -28
rect 11604 -30 11610 22
rect 11958 20 14440 21
rect 14756 20 15006 28
rect 11958 -23 15006 20
rect 11906 -33 11958 -27
rect 14756 -32 15006 -23
rect 15006 -38 15066 -32
rect 12572 -76 12624 -70
rect 8683 -118 12572 -86
rect 6424 -964 6430 -912
rect 6482 -964 6488 -912
rect 7659 -936 7665 -884
rect 7717 -936 7723 -884
rect 8683 -924 8715 -118
rect 12572 -134 12624 -128
rect 13566 -180 13572 -129
rect 13538 -181 13572 -180
rect 13624 -181 13630 -129
rect 13538 -191 13619 -181
rect 9690 -232 13619 -191
rect 9690 -915 9731 -232
rect 14570 -290 14622 -284
rect 10696 -335 14570 -297
rect 9685 -921 9737 -915
rect 8667 -976 8673 -924
rect 8725 -976 8731 -924
rect 10696 -924 10734 -335
rect 14570 -348 14622 -342
rect 15581 -435 15587 -428
rect 11695 -473 15587 -435
rect 11695 -924 11733 -473
rect 15581 -480 15587 -473
rect 15639 -480 15645 -428
rect 16594 -544 16646 -538
rect 12712 -589 16594 -551
rect 12712 -908 12750 -589
rect 16594 -602 16646 -596
rect 17597 -704 17603 -698
rect 13714 -744 17603 -704
rect 9685 -979 9737 -973
rect 10683 -976 10689 -924
rect 10741 -976 10747 -924
rect 11688 -930 11740 -924
rect 12699 -960 12705 -908
rect 12757 -960 12763 -908
rect 13714 -928 13754 -744
rect 17597 -750 17603 -744
rect 17655 -750 17661 -698
rect 18606 -858 18646 527
rect 14727 -898 18646 -858
rect 13708 -934 13760 -928
rect 11688 -988 11740 -982
rect 13708 -992 13760 -986
rect 326 -1088 388 -1076
rect 14727 -1077 14767 -898
rect 326 -1095 332 -1088
rect 319 -1147 325 -1095
rect 326 -1154 332 -1147
rect 382 -1154 388 -1088
rect 3756 -1086 3846 -1082
rect 3756 -1088 3782 -1086
rect 3756 -1140 3768 -1088
rect 3835 -1139 3846 -1086
rect 14702 -1083 14792 -1077
rect 14702 -1123 14714 -1083
rect 14780 -1123 14792 -1083
rect 8090 -1130 8168 -1124
rect 14702 -1129 14792 -1123
rect 3834 -1140 3846 -1139
rect 3756 -1146 3846 -1140
rect 326 -1166 388 -1154
rect 8084 -1182 8090 -1130
rect 8168 -1182 8174 -1130
rect 11120 -1150 11126 -1130
rect 9098 -1155 9176 -1150
rect 10106 -1153 10184 -1150
rect 8084 -1183 8174 -1182
rect 9092 -1156 9182 -1155
rect 8090 -1188 8168 -1183
rect 9092 -1208 9098 -1156
rect 9176 -1208 9182 -1156
rect 10100 -1156 10190 -1153
rect 11114 -1156 11126 -1150
rect 10100 -1208 10106 -1156
rect 10184 -1208 10190 -1156
rect 11108 -1208 11114 -1156
rect 11186 -1156 11192 -1130
rect 11192 -1208 11198 -1156
rect 12133 -1189 12139 -1137
rect 12191 -1189 12197 -1137
rect 13136 -1198 13142 -1146
rect 13194 -1198 13200 -1146
rect 14136 -1189 14142 -1137
rect 14194 -1189 14200 -1137
rect 15166 -1188 15172 -1136
rect 15224 -1188 15230 -1136
rect 36 -1218 126 -1212
rect 36 -1284 48 -1218
rect 114 -1284 126 -1218
rect 36 -1289 55 -1284
rect 107 -1289 126 -1284
rect 36 -1290 126 -1289
rect 3494 -1218 3572 -1212
rect 9098 -1214 9176 -1208
rect 10106 -1214 10184 -1208
rect 11114 -1214 11192 -1208
rect 3494 -1284 3500 -1218
rect 3566 -1284 3572 -1218
rect 7221 -1282 7227 -1230
rect 7279 -1282 7285 -1230
rect 7652 -1282 7730 -1276
rect 8223 -1280 8229 -1228
rect 8281 -1280 8287 -1228
rect 8660 -1259 8738 -1253
rect 3494 -1290 3572 -1284
rect 2958 -1404 3048 -1398
rect 2958 -1457 2970 -1404
rect 3036 -1457 3048 -1404
rect 3294 -1400 3384 -1394
rect 3294 -1405 3306 -1400
rect 3372 -1405 3384 -1400
rect 3294 -1457 3300 -1405
rect 3378 -1457 3384 -1405
rect 2958 -1463 3048 -1457
rect 3300 -1463 3378 -1457
rect 2977 -1517 3030 -1463
rect 2972 -1570 2978 -1517
rect 3030 -1570 3036 -1517
rect 2977 -1603 3030 -1570
rect 64 -1656 3030 -1603
rect 3508 -1614 3557 -1290
rect 7646 -1334 7652 -1282
rect 7730 -1334 7736 -1282
rect 8654 -1311 8660 -1259
rect 8738 -1311 8744 -1259
rect 9235 -1278 9241 -1226
rect 9293 -1278 9299 -1226
rect 9680 -1299 9686 -1247
rect 9738 -1299 9744 -1247
rect 10248 -1280 10254 -1228
rect 10306 -1280 10312 -1228
rect 10676 -1250 10754 -1244
rect 10670 -1301 10676 -1251
rect 10754 -1301 10760 -1251
rect 11254 -1276 11260 -1224
rect 11312 -1276 11318 -1224
rect 11682 -1300 11688 -1248
rect 11740 -1300 11746 -1248
rect 12269 -1278 12275 -1226
rect 12327 -1278 12333 -1226
rect 12692 -1262 12770 -1256
rect 10676 -1308 10754 -1302
rect 8654 -1312 8744 -1311
rect 8660 -1317 8738 -1312
rect 12686 -1313 12692 -1263
rect 12770 -1313 12776 -1263
rect 13268 -1274 13274 -1222
rect 13326 -1274 13332 -1222
rect 13702 -1288 13708 -1236
rect 13760 -1288 13766 -1236
rect 14283 -1280 14289 -1228
rect 14341 -1280 14347 -1228
rect 12692 -1320 12770 -1314
rect 7646 -1336 7658 -1334
rect 7724 -1336 7736 -1334
rect 7646 -1342 7736 -1336
rect 6746 -1406 6836 -1400
rect 6410 -1416 6500 -1410
rect 6410 -1421 6422 -1416
rect 6488 -1421 6500 -1416
rect 6410 -1473 6416 -1421
rect 6494 -1473 6500 -1421
rect 6746 -1412 6758 -1406
rect 6824 -1412 6836 -1406
rect 6746 -1465 6752 -1412
rect 6830 -1465 6836 -1412
rect 6752 -1471 6830 -1465
rect 6416 -1479 6494 -1473
rect 5602 -1554 5608 -1502
rect 5664 -1503 5670 -1502
rect 9335 -1503 9341 -1499
rect 5664 -1508 6386 -1503
rect 6524 -1508 9341 -1503
rect 5664 -1546 9341 -1508
rect 5664 -1554 5670 -1546
rect 9335 -1551 9341 -1546
rect 9393 -1551 9399 -1499
rect 15159 -1602 15211 -1596
rect 64 -1978 117 -1656
rect 3508 -1663 6480 -1614
rect 6880 -1656 6886 -1604
rect 6938 -1612 6944 -1604
rect 9106 -1612 9112 -1604
rect 6938 -1648 9112 -1612
rect 6938 -1656 6944 -1648
rect 9106 -1656 9112 -1648
rect 9164 -1656 9170 -1604
rect 15159 -1660 15211 -1654
rect 2977 -1760 3448 -1708
rect 3500 -1760 3554 -1708
rect 2977 -1805 3029 -1760
rect 2958 -1811 3048 -1805
rect 3300 -1811 3378 -1805
rect 2958 -1877 2970 -1811
rect 3036 -1877 3048 -1811
rect 3294 -1863 3300 -1811
rect 3378 -1863 3384 -1811
rect 3294 -1864 3306 -1863
rect 3372 -1864 3384 -1863
rect 3294 -1870 3384 -1864
rect 2958 -1883 3048 -1877
rect 3502 -1972 3554 -1760
rect 6431 -1809 6480 -1663
rect 7540 -1757 7592 -1751
rect 10796 -1759 10802 -1756
rect 7592 -1806 10802 -1759
rect 10796 -1808 10802 -1806
rect 10854 -1808 10860 -1756
rect 6410 -1810 6500 -1809
rect 6410 -1815 6430 -1810
rect 6482 -1815 6500 -1810
rect 6752 -1815 6830 -1809
rect 7540 -1815 7592 -1809
rect 6410 -1864 6422 -1815
rect 6488 -1864 6500 -1815
rect 6410 -1870 6500 -1864
rect 6746 -1867 6752 -1815
rect 6830 -1867 6836 -1815
rect 6746 -1872 6758 -1867
rect 6824 -1872 6836 -1867
rect 6746 -1878 6836 -1872
rect 6940 -1899 7030 -1893
rect 6940 -1933 6952 -1899
rect 7018 -1933 7030 -1899
rect 6940 -1939 7030 -1933
rect 9668 -1939 9746 -1933
rect 3494 -1978 3571 -1972
rect 42 -1984 120 -1978
rect 42 -2050 48 -1984
rect 114 -2050 120 -1984
rect 42 -2056 120 -2050
rect 3488 -1984 3578 -1978
rect 3488 -2050 3500 -1984
rect 3566 -2050 3578 -1984
rect 6971 -2041 6999 -1939
rect 7214 -1978 7292 -1972
rect 7652 -1973 7730 -1967
rect 8660 -1973 8738 -1967
rect 7208 -2030 7214 -1978
rect 7292 -2030 7298 -1978
rect 7208 -2034 7220 -2030
rect 7286 -2034 7298 -2030
rect 7646 -2025 7652 -1973
rect 7730 -2025 7736 -1973
rect 7646 -2028 7658 -2025
rect 7724 -2028 7736 -2025
rect 7646 -2034 7736 -2028
rect 7208 -2040 7298 -2034
rect 3488 -2056 3578 -2050
rect 3494 -2062 3571 -2056
rect 310 -2114 388 -2102
rect 310 -2180 316 -2114
rect 382 -2180 388 -2114
rect 310 -2192 388 -2180
rect 3768 -2114 3840 -2102
rect 3768 -2180 3774 -2114
rect 3834 -2180 3840 -2114
rect 3768 -2192 3840 -2180
rect 3608 -2354 3660 -2348
rect 3608 -2412 3660 -2406
rect 3616 -2512 3651 -2412
rect 3783 -2452 3834 -2192
rect 6760 -2289 6766 -2237
rect 6818 -2289 6824 -2237
rect 6767 -2452 6818 -2289
rect 3783 -2503 6818 -2452
rect 6963 -2486 7006 -2041
rect 8226 -2047 8232 -1995
rect 8284 -2047 8290 -1995
rect 8654 -2025 8660 -1973
rect 8738 -2025 8744 -1973
rect 9662 -1991 9668 -1939
rect 9746 -1991 9752 -1939
rect 11684 -1957 11762 -1951
rect 12692 -1955 12770 -1949
rect 10676 -1963 10754 -1957
rect 9662 -1992 9752 -1991
rect 8654 -2041 8666 -2025
rect 8732 -2041 8744 -2025
rect 8654 -2047 8744 -2041
rect 9234 -2044 9240 -1992
rect 9292 -2044 9298 -1992
rect 9668 -1997 9746 -1992
rect 10240 -2041 10246 -1989
rect 10298 -2041 10304 -1989
rect 10670 -2015 10676 -1963
rect 10754 -2015 10760 -1963
rect 10670 -2019 10760 -2015
rect 10676 -2021 10754 -2019
rect 11246 -2048 11252 -1996
rect 11304 -2048 11310 -1996
rect 11678 -2009 11684 -1957
rect 11762 -2009 11768 -1957
rect 11678 -2013 11768 -2009
rect 11684 -2015 11762 -2013
rect 12256 -2039 12262 -1987
rect 12314 -2039 12320 -1987
rect 12686 -2006 12692 -1957
rect 12770 -2006 12776 -1957
rect 13700 -1961 13778 -1955
rect 12692 -2013 12770 -2007
rect 13262 -2046 13268 -1994
rect 13320 -2046 13326 -1994
rect 13694 -2013 13700 -1961
rect 13778 -2013 13784 -1961
rect 14708 -1967 14786 -1961
rect 13700 -2019 13778 -2013
rect 14274 -2039 14280 -1987
rect 14332 -2039 14338 -1987
rect 14702 -2019 14708 -1967
rect 14786 -2019 14792 -1967
rect 14702 -2024 14792 -2019
rect 14708 -2025 14786 -2024
rect 15165 -2060 15205 -1660
rect 8108 -2128 8114 -2076
rect 8166 -2128 8172 -2076
rect 9098 -2128 9104 -2076
rect 9156 -2128 9162 -2076
rect 10108 -2124 10114 -2072
rect 10166 -2124 10172 -2072
rect 11132 -2073 11184 -2067
rect 14151 -2069 14203 -2063
rect 11132 -2131 11184 -2125
rect 12134 -2126 12140 -2074
rect 12192 -2126 12198 -2074
rect 13144 -2082 13196 -2076
rect 15140 -2066 15230 -2060
rect 15140 -2106 15152 -2066
rect 15218 -2106 15230 -2066
rect 15140 -2112 15230 -2106
rect 14151 -2127 14203 -2121
rect 13144 -2140 13196 -2134
rect 7108 -2185 7160 -2179
rect 7326 -2185 7332 -2184
rect 7160 -2236 7332 -2185
rect 7384 -2236 7390 -2184
rect 7108 -2243 7160 -2237
rect 7090 -2349 7150 -2343
rect 7150 -2405 8114 -2353
rect 8166 -2405 8172 -2353
rect 7090 -2415 7150 -2409
rect 15313 -2483 15365 -2477
rect -27 -2547 3651 -2512
rect 6963 -2529 15313 -2486
rect 7296 -2531 15313 -2529
rect 15313 -2541 15365 -2535
<< via1 >>
rect 308 580 316 632
rect 316 580 360 632
rect 10217 940 10269 992
rect 3781 580 3833 632
rect 11542 571 11620 572
rect 11542 526 11548 571
rect 11548 526 11614 571
rect 11614 526 11620 571
rect 11542 520 11620 526
rect 12572 584 12624 590
rect 12572 544 12578 584
rect 12578 544 12618 584
rect 12618 544 12624 584
rect 12572 538 12624 544
rect 13558 567 13636 572
rect 13558 526 13564 567
rect 13564 526 13630 567
rect 13630 526 13636 567
rect 13558 520 13636 526
rect 14570 580 14622 586
rect 14570 540 14576 580
rect 14576 540 14616 580
rect 14616 540 14622 580
rect 14570 534 14622 540
rect 15574 564 15652 571
rect 15574 526 15580 564
rect 15580 526 15646 564
rect 15646 526 15652 564
rect 15574 519 15652 526
rect 16594 580 16646 586
rect 16594 540 16600 580
rect 16600 540 16640 580
rect 16640 540 16646 580
rect 16594 534 16646 540
rect 17590 566 17668 572
rect 17590 526 17596 566
rect 17596 526 17662 566
rect 17662 526 17668 566
rect 17590 520 17668 526
rect 6970 444 7018 494
rect 7018 444 7022 494
rect 6970 442 7022 444
rect 10688 498 10740 504
rect 10688 458 10694 498
rect 10694 458 10734 498
rect 10734 458 10740 498
rect 10688 452 10740 458
rect 11680 499 11732 505
rect 11680 459 11686 499
rect 11686 459 11726 499
rect 11726 459 11732 499
rect 11680 453 11732 459
rect 12690 501 12742 507
rect 12690 461 12696 501
rect 12696 461 12736 501
rect 12736 461 12742 501
rect 12690 455 12742 461
rect 13694 501 13746 507
rect 13694 461 13700 501
rect 13700 461 13740 501
rect 13740 461 13746 501
rect 13694 455 13746 461
rect 14708 497 14760 503
rect 14708 457 14714 497
rect 14714 457 14754 497
rect 14754 457 14760 497
rect 14708 451 14760 457
rect 15714 499 15766 505
rect 15714 459 15720 499
rect 15720 459 15760 499
rect 15760 459 15766 499
rect 15714 453 15766 459
rect 16720 503 16772 509
rect 16720 463 16726 503
rect 16726 463 16766 503
rect 16766 463 16772 503
rect 16720 457 16772 463
rect 17730 497 17782 503
rect 17730 457 17736 497
rect 17736 457 17776 497
rect 17776 457 17782 497
rect 17730 451 17782 457
rect -35 329 17 381
rect 3300 311 3378 320
rect 3300 277 3306 311
rect 3306 277 3372 311
rect 3372 277 3378 311
rect 3300 268 3378 277
rect 2977 128 3029 180
rect 6416 277 6422 323
rect 6422 277 6488 323
rect 6488 277 6494 323
rect 6416 271 6494 277
rect 6752 265 6758 311
rect 6758 265 6824 311
rect 6824 265 6830 311
rect 6752 259 6830 265
rect 9868 308 9946 311
rect 9868 265 9874 308
rect 9874 265 9940 308
rect 9940 265 9946 308
rect 9868 259 9946 265
rect 10204 326 10282 332
rect 10204 280 10210 326
rect 10210 280 10276 326
rect 10276 280 10282 326
rect 2964 -89 3042 -83
rect 2964 -130 2970 -89
rect 2970 -130 3036 -89
rect 3036 -130 3042 -89
rect 2964 -135 3042 -130
rect 3300 -87 3378 -81
rect 3300 -133 3306 -87
rect 3306 -133 3372 -87
rect 3372 -133 3378 -87
rect 6752 -133 6758 -87
rect 6758 -133 6824 -87
rect 6824 -133 6830 -87
rect 6752 -139 6830 -133
rect 6951 -190 7003 -138
rect 327 -445 379 -393
rect 3782 -440 3834 -388
rect 3676 -658 3728 -606
rect 3890 -657 3942 -605
rect 6650 -656 6702 -604
rect 6870 -789 6922 -737
rect 11552 -30 11604 22
rect 11906 -27 11958 25
rect 15006 -32 15066 28
rect 6430 -964 6482 -912
rect 7665 -936 7717 -884
rect 12572 -128 12624 -76
rect 13572 -181 13624 -129
rect 8673 -976 8725 -924
rect 9685 -973 9737 -921
rect 14570 -342 14622 -290
rect 15587 -480 15639 -428
rect 16594 -596 16646 -544
rect 10689 -976 10741 -924
rect 11688 -982 11740 -930
rect 12705 -960 12757 -908
rect 17603 -750 17655 -698
rect 13708 -986 13760 -934
rect 325 -1147 332 -1095
rect 332 -1147 377 -1095
rect 3782 -1088 3835 -1086
rect 3782 -1139 3834 -1088
rect 3834 -1139 3835 -1088
rect 8090 -1136 8168 -1130
rect 8090 -1177 8096 -1136
rect 8096 -1177 8162 -1136
rect 8162 -1177 8168 -1136
rect 8090 -1182 8168 -1177
rect 11126 -1150 11186 -1130
rect 9098 -1161 9176 -1156
rect 9098 -1202 9104 -1161
rect 9104 -1202 9170 -1161
rect 9170 -1202 9176 -1161
rect 9098 -1208 9176 -1202
rect 11126 -1156 11132 -1150
rect 10106 -1159 10184 -1156
rect 10106 -1202 10112 -1159
rect 10112 -1202 10178 -1159
rect 10178 -1202 10184 -1159
rect 10106 -1208 10184 -1202
rect 11114 -1162 11132 -1156
rect 11132 -1162 11180 -1150
rect 11180 -1156 11186 -1150
rect 11180 -1162 11192 -1156
rect 11114 -1202 11120 -1162
rect 11120 -1202 11186 -1162
rect 11186 -1202 11192 -1162
rect 11114 -1208 11192 -1202
rect 12139 -1143 12191 -1137
rect 12139 -1183 12145 -1143
rect 12145 -1183 12185 -1143
rect 12185 -1183 12191 -1143
rect 12139 -1189 12191 -1183
rect 13142 -1152 13194 -1146
rect 13142 -1192 13148 -1152
rect 13148 -1192 13188 -1152
rect 13188 -1192 13194 -1152
rect 13142 -1198 13194 -1192
rect 14142 -1143 14194 -1137
rect 14142 -1183 14148 -1143
rect 14148 -1183 14188 -1143
rect 14188 -1183 14194 -1143
rect 14142 -1189 14194 -1183
rect 15172 -1142 15224 -1136
rect 15172 -1182 15178 -1142
rect 15178 -1182 15218 -1142
rect 15218 -1182 15224 -1142
rect 15172 -1188 15224 -1182
rect 55 -1284 107 -1237
rect 55 -1289 107 -1284
rect 7227 -1236 7279 -1230
rect 7227 -1276 7233 -1236
rect 7233 -1276 7273 -1236
rect 7273 -1276 7279 -1236
rect 7227 -1282 7279 -1276
rect 8229 -1234 8281 -1228
rect 8229 -1274 8235 -1234
rect 8235 -1274 8275 -1234
rect 8275 -1274 8281 -1234
rect 8229 -1280 8281 -1274
rect 3300 -1451 3306 -1405
rect 3306 -1451 3372 -1405
rect 3372 -1451 3378 -1405
rect 3300 -1457 3378 -1451
rect 2978 -1570 3030 -1517
rect 7652 -1288 7730 -1282
rect 7652 -1334 7658 -1288
rect 7658 -1334 7724 -1288
rect 7724 -1334 7730 -1288
rect 8660 -1265 8738 -1259
rect 8660 -1306 8666 -1265
rect 8666 -1306 8732 -1265
rect 8732 -1306 8738 -1265
rect 8660 -1311 8738 -1306
rect 9241 -1232 9293 -1226
rect 9241 -1272 9247 -1232
rect 9247 -1272 9287 -1232
rect 9287 -1272 9293 -1232
rect 9241 -1278 9293 -1272
rect 9686 -1253 9738 -1247
rect 9686 -1293 9692 -1253
rect 9692 -1293 9732 -1253
rect 9732 -1293 9738 -1253
rect 9686 -1299 9738 -1293
rect 10254 -1234 10306 -1228
rect 10254 -1274 10260 -1234
rect 10260 -1274 10300 -1234
rect 10300 -1274 10306 -1234
rect 10254 -1280 10306 -1274
rect 10676 -1257 10754 -1250
rect 10676 -1295 10682 -1257
rect 10682 -1295 10748 -1257
rect 10748 -1295 10754 -1257
rect 10676 -1302 10754 -1295
rect 11260 -1230 11312 -1224
rect 11260 -1270 11266 -1230
rect 11266 -1270 11306 -1230
rect 11306 -1270 11312 -1230
rect 11260 -1276 11312 -1270
rect 11688 -1254 11740 -1248
rect 11688 -1294 11700 -1254
rect 11700 -1294 11734 -1254
rect 11734 -1294 11740 -1254
rect 11688 -1300 11740 -1294
rect 12275 -1232 12327 -1226
rect 12275 -1272 12281 -1232
rect 12281 -1272 12321 -1232
rect 12321 -1272 12327 -1232
rect 12275 -1278 12327 -1272
rect 12692 -1269 12770 -1262
rect 12692 -1307 12698 -1269
rect 12698 -1307 12764 -1269
rect 12764 -1307 12770 -1269
rect 12692 -1314 12770 -1307
rect 13274 -1228 13326 -1222
rect 13274 -1268 13280 -1228
rect 13280 -1268 13320 -1228
rect 13320 -1268 13326 -1228
rect 13274 -1274 13326 -1268
rect 13708 -1242 13760 -1236
rect 13708 -1282 13714 -1242
rect 13714 -1282 13754 -1242
rect 13754 -1282 13760 -1242
rect 13708 -1288 13760 -1282
rect 14289 -1234 14341 -1228
rect 14289 -1274 14295 -1234
rect 14295 -1274 14335 -1234
rect 14335 -1274 14341 -1234
rect 14289 -1280 14341 -1274
rect 6416 -1467 6422 -1421
rect 6422 -1467 6488 -1421
rect 6488 -1467 6494 -1421
rect 6416 -1473 6494 -1467
rect 6752 -1459 6758 -1412
rect 6758 -1459 6824 -1412
rect 6824 -1459 6830 -1412
rect 6752 -1465 6830 -1459
rect 5608 -1554 5664 -1502
rect 9341 -1551 9393 -1499
rect 6886 -1656 6938 -1604
rect 9112 -1656 9164 -1604
rect 15159 -1654 15211 -1602
rect 3448 -1760 3500 -1708
rect 3300 -1817 3378 -1811
rect 3300 -1863 3306 -1817
rect 3306 -1863 3372 -1817
rect 3372 -1863 3378 -1817
rect 7540 -1809 7592 -1757
rect 10802 -1808 10854 -1756
rect 6430 -1815 6482 -1810
rect 6430 -1862 6482 -1815
rect 6752 -1821 6830 -1815
rect 6752 -1867 6758 -1821
rect 6758 -1867 6824 -1821
rect 6824 -1867 6830 -1821
rect 7214 -1984 7292 -1978
rect 7214 -2030 7220 -1984
rect 7220 -2030 7286 -1984
rect 7286 -2030 7292 -1984
rect 7652 -1979 7730 -1973
rect 7652 -2025 7658 -1979
rect 7658 -2025 7724 -1979
rect 7724 -2025 7730 -1979
rect 329 -2175 381 -2123
rect 3608 -2406 3660 -2354
rect 6766 -2289 6818 -2237
rect 8232 -2001 8284 -1995
rect 8232 -2041 8238 -2001
rect 8238 -2041 8278 -2001
rect 8278 -2041 8284 -2001
rect 8232 -2047 8284 -2041
rect 8660 -1979 8738 -1973
rect 8660 -2025 8666 -1979
rect 8666 -2025 8732 -1979
rect 8732 -2025 8738 -1979
rect 9668 -1945 9746 -1939
rect 9668 -1986 9674 -1945
rect 9674 -1986 9740 -1945
rect 9740 -1986 9746 -1945
rect 9668 -1991 9746 -1986
rect 9240 -1998 9292 -1992
rect 9240 -2038 9246 -1998
rect 9246 -2038 9286 -1998
rect 9286 -2038 9292 -1998
rect 9240 -2044 9292 -2038
rect 10246 -1995 10298 -1989
rect 10246 -2035 10252 -1995
rect 10252 -2035 10292 -1995
rect 10292 -2035 10298 -1995
rect 10246 -2041 10298 -2035
rect 10676 -1969 10754 -1963
rect 10676 -2013 10682 -1969
rect 10682 -2013 10748 -1969
rect 10748 -2013 10754 -1969
rect 10676 -2015 10754 -2013
rect 11252 -2002 11304 -1996
rect 11252 -2042 11258 -2002
rect 11258 -2042 11298 -2002
rect 11298 -2042 11304 -2002
rect 11252 -2048 11304 -2042
rect 11684 -1963 11762 -1957
rect 11684 -2007 11690 -1963
rect 11690 -2007 11756 -1963
rect 11756 -2007 11762 -1963
rect 11684 -2009 11762 -2007
rect 12262 -1993 12314 -1987
rect 12262 -2033 12268 -1993
rect 12268 -2033 12308 -1993
rect 12308 -2033 12314 -1993
rect 12262 -2039 12314 -2033
rect 12692 -1963 12770 -1955
rect 12692 -2000 12698 -1963
rect 12698 -2000 12764 -1963
rect 12764 -2000 12770 -1963
rect 12692 -2007 12770 -2000
rect 13268 -2000 13320 -1994
rect 13268 -2040 13274 -2000
rect 13274 -2040 13314 -2000
rect 13314 -2040 13320 -2000
rect 13268 -2046 13320 -2040
rect 13700 -1967 13778 -1961
rect 13700 -2007 13706 -1967
rect 13706 -2007 13772 -1967
rect 13772 -2007 13778 -1967
rect 13700 -2013 13778 -2007
rect 14280 -1993 14332 -1987
rect 14280 -2033 14286 -1993
rect 14286 -2033 14326 -1993
rect 14326 -2033 14332 -1993
rect 14280 -2039 14332 -2033
rect 14708 -1973 14786 -1967
rect 14708 -2018 14714 -1973
rect 14714 -2018 14780 -1973
rect 14780 -2018 14786 -1973
rect 14708 -2019 14786 -2018
rect 8114 -2082 8166 -2076
rect 8114 -2122 8120 -2082
rect 8120 -2122 8160 -2082
rect 8160 -2122 8166 -2082
rect 8114 -2128 8166 -2122
rect 9104 -2082 9156 -2076
rect 9104 -2122 9110 -2082
rect 9110 -2122 9150 -2082
rect 9150 -2122 9156 -2082
rect 9104 -2128 9156 -2122
rect 10114 -2078 10166 -2072
rect 10114 -2118 10120 -2078
rect 10120 -2118 10160 -2078
rect 10160 -2118 10166 -2078
rect 10114 -2124 10166 -2118
rect 11132 -2079 11184 -2073
rect 11132 -2119 11138 -2079
rect 11138 -2119 11178 -2079
rect 11178 -2119 11184 -2079
rect 11132 -2125 11184 -2119
rect 12140 -2080 12192 -2074
rect 12140 -2120 12146 -2080
rect 12146 -2120 12186 -2080
rect 12186 -2120 12192 -2080
rect 12140 -2126 12192 -2120
rect 14151 -2075 14203 -2069
rect 13144 -2088 13196 -2082
rect 13144 -2128 13150 -2088
rect 13150 -2128 13190 -2088
rect 13190 -2128 13196 -2088
rect 14151 -2115 14157 -2075
rect 14157 -2115 14197 -2075
rect 14197 -2115 14203 -2075
rect 14151 -2121 14203 -2115
rect 13144 -2134 13196 -2128
rect 7108 -2237 7160 -2185
rect 7332 -2236 7384 -2184
rect 7090 -2409 7150 -2349
rect 8114 -2405 8166 -2353
rect 15313 -2535 15365 -2483
<< metal2 >>
rect 10217 992 10269 998
rect 10269 940 10304 942
rect 10217 934 10304 940
rect 10218 911 10304 934
rect 10218 861 18741 911
rect 308 632 360 638
rect 308 574 360 580
rect 3781 632 3833 638
rect 3781 574 3833 580
rect -35 381 17 387
rect 320 373 348 574
rect 17 338 349 373
rect -35 323 17 329
rect 320 308 348 338
rect 3294 308 3300 320
rect 320 280 3300 308
rect 3294 268 3300 280
rect 3378 268 3384 320
rect -11 175 2911 215
rect 2971 175 2977 180
rect -11 173 2977 175
rect -11 -1135 31 173
rect 2869 133 2977 173
rect 2971 128 2977 133
rect 3029 128 3042 180
rect 3782 115 3831 574
rect 6964 492 6970 494
rect 6431 443 6970 492
rect 6431 323 6480 443
rect 6410 271 6416 323
rect 6494 271 6500 323
rect 6746 259 6752 311
rect 6830 259 6836 311
rect 6767 115 6816 259
rect 314 40 323 100
rect 383 95 392 100
rect 383 44 3365 95
rect 3782 66 6816 115
rect 6877 115 6926 443
rect 6964 442 6970 443
rect 7022 442 7028 494
rect 10218 332 10268 861
rect 10692 718 17777 761
rect 10692 510 10735 718
rect 11536 520 11542 572
rect 11620 520 11626 572
rect 10688 504 10740 510
rect 10688 446 10740 452
rect 9862 259 9868 311
rect 9946 259 9952 311
rect 10198 280 10204 332
rect 10282 280 10288 332
rect 9886 154 9929 259
rect 10692 154 10735 446
rect 6877 66 9728 115
rect 9886 111 10735 154
rect 383 40 392 44
rect 327 -387 378 40
rect 3314 -81 3365 44
rect 6746 18 6794 66
rect 7135 18 7144 22
rect 6746 -30 7144 18
rect 7135 -34 7144 -30
rect 7200 -34 7209 22
rect 2958 -135 2964 -83
rect 3042 -135 3048 -83
rect 3294 -133 3300 -81
rect 3378 -133 3384 -81
rect 327 -393 379 -387
rect 327 -451 379 -445
rect 2983 -693 3024 -135
rect 6746 -139 6752 -87
rect 6830 -139 6836 -87
rect 6766 -140 6836 -139
rect 6951 -138 7003 -132
rect 3782 -388 3834 -382
rect 3782 -446 3834 -440
rect 6766 -419 6816 -140
rect 7003 -189 9451 -139
rect 6951 -196 7003 -190
rect 9149 -419 9158 -414
rect 3676 -606 3728 -600
rect 3676 -664 3728 -658
rect 3681 -693 3722 -664
rect -41 -1177 31 -1135
rect 60 -734 3722 -693
rect -41 -1353 1 -1177
rect 60 -1231 101 -734
rect 3783 -751 3833 -446
rect 6766 -469 9158 -419
rect 3890 -605 3942 -599
rect 6644 -610 6650 -604
rect 3942 -651 6650 -610
rect 6644 -656 6650 -651
rect 6702 -656 6708 -604
rect 3890 -663 3942 -657
rect 6766 -751 6816 -469
rect 9149 -474 9158 -469
rect 9218 -474 9227 -414
rect 3783 -801 6816 -751
rect 6870 -737 6922 -731
rect 6922 -783 8150 -742
rect 6870 -795 6922 -789
rect 325 -825 3365 -821
rect 325 -834 3370 -825
rect 325 -872 3310 -834
rect 325 -1089 376 -872
rect 7665 -884 7717 -878
rect 3310 -903 3370 -894
rect 6909 -898 6918 -894
rect 325 -1095 377 -1089
rect 325 -1153 377 -1147
rect 55 -1237 107 -1231
rect 55 -1295 107 -1289
rect -41 -1399 33 -1353
rect -17 -2461 33 -1399
rect 3314 -1405 3365 -903
rect 6765 -904 6918 -898
rect 6433 -906 6918 -904
rect 6430 -912 6918 -906
rect 6482 -946 6918 -912
rect 6765 -951 6918 -946
rect 6765 -952 6818 -951
rect 6909 -954 6918 -951
rect 6978 -954 6987 -894
rect 7665 -942 7717 -936
rect 6430 -970 6482 -964
rect 3782 -1086 3835 -1080
rect 3294 -1457 3300 -1405
rect 3378 -1457 3384 -1405
rect 2978 -1517 3030 -1511
rect 3347 -1524 3356 -1513
rect 3030 -1562 3356 -1524
rect 2978 -1576 3030 -1570
rect 3347 -1573 3356 -1562
rect 3416 -1573 3425 -1513
rect 3782 -1605 3835 -1139
rect 6430 -1421 6481 -970
rect 7227 -1230 7279 -1224
rect 7667 -1282 7715 -942
rect 8109 -1130 8150 -783
rect 9401 -749 9451 -189
rect 9679 -601 9728 66
rect 10218 -431 10268 111
rect 11559 28 11604 520
rect 11684 511 11727 718
rect 12572 590 12624 596
rect 12572 532 12624 538
rect 11680 505 11732 511
rect 11680 447 11732 453
rect 11552 22 11604 28
rect 11900 -27 11906 25
rect 11958 -27 11964 25
rect 11552 -36 11604 -30
rect 10359 -144 10368 -84
rect 10428 -92 10437 -84
rect 11910 -92 11954 -27
rect 12582 -76 12614 532
rect 12694 513 12737 718
rect 13552 520 13558 572
rect 13636 520 13642 572
rect 12690 507 12742 513
rect 12690 449 12742 455
rect 10428 -136 11954 -92
rect 12566 -128 12572 -76
rect 12624 -128 12630 -76
rect 13577 -123 13618 520
rect 13698 513 13741 718
rect 14570 586 14622 592
rect 14570 528 14622 534
rect 13694 507 13746 513
rect 13694 449 13746 455
rect 13572 -129 13624 -123
rect 10428 -144 10437 -136
rect 13572 -187 13624 -181
rect 14577 -290 14615 528
rect 14712 509 14755 718
rect 15568 519 15574 571
rect 15652 519 15658 571
rect 14708 503 14760 509
rect 14708 445 14760 451
rect 15008 28 15064 35
rect 15000 -32 15006 28
rect 15066 -32 15072 28
rect 15008 -39 15064 -32
rect 14564 -342 14570 -290
rect 14622 -342 14628 -290
rect 15594 -422 15632 519
rect 15718 511 15761 718
rect 16594 586 16646 592
rect 16594 528 16646 534
rect 15714 505 15766 511
rect 15714 447 15766 453
rect 15587 -428 15639 -422
rect 10218 -481 15223 -431
rect 9679 -650 14192 -601
rect 14886 -604 14946 -602
rect 9401 -799 13193 -749
rect 12136 -896 12192 -887
rect 8673 -924 8725 -918
rect 9679 -973 9685 -921
rect 9737 -973 9743 -921
rect 10689 -924 10741 -918
rect 8673 -982 8725 -976
rect 8084 -1182 8090 -1130
rect 8168 -1182 8174 -1130
rect 7227 -1288 7279 -1282
rect 6626 -1344 6930 -1308
rect 5444 -1468 5782 -1432
rect 3913 -1540 3922 -1484
rect 3978 -1494 3987 -1484
rect 5444 -1494 5480 -1468
rect 3978 -1530 5480 -1494
rect 5608 -1502 5664 -1496
rect 3978 -1540 3987 -1530
rect 5599 -1558 5608 -1502
rect 5664 -1558 5673 -1502
rect 5746 -1508 5782 -1468
rect 6410 -1473 6416 -1421
rect 6494 -1473 6500 -1421
rect 6626 -1508 6662 -1344
rect 6765 -1412 6818 -1400
rect 6746 -1465 6752 -1412
rect 6830 -1465 6836 -1412
rect 5746 -1544 6662 -1508
rect 5608 -1560 5664 -1558
rect 5905 -1605 5958 -1604
rect 6765 -1605 6818 -1465
rect 6894 -1598 6930 -1344
rect 331 -1660 3363 -1613
rect 3782 -1658 6818 -1605
rect 6886 -1604 6938 -1598
rect 331 -2117 378 -1660
rect 3316 -1811 3363 -1660
rect 5905 -1698 5958 -1658
rect 6886 -1662 6938 -1656
rect 7228 -1636 7277 -1288
rect 7646 -1334 7652 -1282
rect 7730 -1334 7736 -1282
rect 7228 -1685 7716 -1636
rect 3448 -1708 3500 -1702
rect 5597 -1708 5606 -1704
rect 3500 -1760 5606 -1708
rect 3448 -1766 3500 -1760
rect 5597 -1764 5606 -1760
rect 5666 -1764 5675 -1704
rect 5902 -1707 5962 -1698
rect 5902 -1776 5962 -1767
rect 6298 -1740 7013 -1693
rect 3294 -1863 3300 -1811
rect 3378 -1863 3384 -1811
rect 3316 -1918 3363 -1863
rect 6298 -1918 6345 -1740
rect 6966 -1760 7013 -1740
rect 7534 -1760 7540 -1757
rect 6418 -1810 6490 -1804
rect 6966 -1807 7540 -1760
rect 6418 -1812 6430 -1810
rect 6482 -1812 6490 -1810
rect 6417 -1868 6426 -1812
rect 6482 -1868 6491 -1812
rect 6762 -1815 6822 -1808
rect 7534 -1809 7540 -1807
rect 7592 -1809 7598 -1757
rect 6746 -1867 6752 -1815
rect 6830 -1867 6836 -1815
rect 3316 -1965 6345 -1918
rect 329 -2123 381 -2117
rect 329 -2181 381 -2175
rect 6766 -2186 6817 -1867
rect 7667 -1973 7716 -1685
rect 8109 -1733 8150 -1182
rect 8229 -1228 8281 -1222
rect 8683 -1259 8715 -982
rect 9092 -1208 9098 -1156
rect 9176 -1208 9182 -1156
rect 8229 -1286 8281 -1280
rect 8232 -1622 8277 -1286
rect 8654 -1311 8660 -1259
rect 8738 -1311 8744 -1259
rect 9117 -1550 9158 -1208
rect 9241 -1226 9293 -1220
rect 9691 -1241 9732 -973
rect 10689 -982 10741 -976
rect 11682 -982 11688 -930
rect 11740 -982 11746 -930
rect 12136 -961 12192 -952
rect 12705 -908 12757 -902
rect 10100 -1208 10106 -1156
rect 10184 -1208 10190 -1156
rect 9241 -1284 9293 -1278
rect 9686 -1247 9738 -1241
rect 9120 -1598 9156 -1550
rect 9112 -1604 9164 -1598
rect 8232 -1667 8722 -1622
rect 9246 -1612 9287 -1284
rect 9686 -1305 9738 -1299
rect 9341 -1499 9393 -1493
rect 10124 -1504 10167 -1208
rect 10254 -1228 10306 -1222
rect 10696 -1250 10734 -982
rect 11126 -1072 11186 -1070
rect 11119 -1128 11128 -1072
rect 11184 -1128 11193 -1072
rect 11126 -1130 11186 -1128
rect 11108 -1208 11114 -1156
rect 11192 -1208 11198 -1156
rect 10254 -1286 10306 -1280
rect 9393 -1547 10167 -1504
rect 9341 -1557 9393 -1551
rect 9246 -1653 9728 -1612
rect 9112 -1662 9164 -1656
rect 8109 -1774 8278 -1733
rect 7208 -2030 7214 -1978
rect 7292 -2030 7298 -1978
rect 7646 -2025 7652 -1973
rect 7730 -2025 7736 -1973
rect 8237 -1989 8278 -1774
rect 8677 -1973 8722 -1667
rect 9120 -1746 9156 -1662
rect 9120 -1782 9284 -1746
rect 8232 -1995 8284 -1989
rect 7102 -2186 7108 -2185
rect 6766 -2237 7108 -2186
rect 7160 -2237 7166 -2185
rect 6766 -2295 6818 -2289
rect 6904 -2349 6960 -2342
rect 3602 -2406 3608 -2354
rect 3660 -2362 3666 -2354
rect 6603 -2362 6612 -2349
rect 3660 -2397 6612 -2362
rect 3660 -2406 3666 -2397
rect 6603 -2409 6612 -2397
rect 6672 -2409 6681 -2349
rect 6902 -2351 7090 -2349
rect 6902 -2407 6904 -2351
rect 6960 -2407 7090 -2351
rect 6902 -2409 7090 -2407
rect 7150 -2409 7156 -2349
rect 6904 -2416 6960 -2409
rect 7228 -2461 7278 -2030
rect 8654 -2025 8660 -1973
rect 8738 -2025 8744 -1973
rect 9248 -1986 9284 -1782
rect 9687 -1939 9728 -1653
rect 10124 -1736 10167 -1547
rect 10258 -1608 10302 -1286
rect 10670 -1302 10676 -1250
rect 10754 -1302 10760 -1250
rect 10258 -1652 10737 -1608
rect 10124 -1779 10293 -1736
rect 10030 -1914 10086 -1905
rect 9240 -1992 9292 -1986
rect 9662 -1991 9668 -1939
rect 9746 -1991 9752 -1939
rect 10086 -1964 10162 -1920
rect 10030 -1979 10086 -1970
rect 8232 -2053 8284 -2047
rect 9240 -2050 9292 -2044
rect 10118 -2066 10162 -1964
rect 10250 -1983 10293 -1779
rect 10693 -1963 10737 -1652
rect 10802 -1756 10854 -1750
rect 10854 -1805 11055 -1758
rect 11133 -1760 11173 -1208
rect 11260 -1224 11312 -1218
rect 11695 -1242 11733 -982
rect 12142 -1131 12187 -961
rect 12705 -966 12757 -960
rect 12139 -1137 12191 -1131
rect 12139 -1195 12191 -1189
rect 11260 -1282 11312 -1276
rect 11688 -1248 11740 -1242
rect 11264 -1606 11308 -1282
rect 11688 -1306 11740 -1300
rect 11264 -1650 11745 -1606
rect 11133 -1800 11298 -1760
rect 10802 -1814 10854 -1808
rect 10246 -1989 10298 -1983
rect 10670 -2015 10676 -1963
rect 10754 -2015 10760 -1963
rect 10246 -2047 10298 -2041
rect 8114 -2076 8166 -2070
rect 7332 -2184 7384 -2178
rect 7943 -2184 7952 -2179
rect 7384 -2235 7952 -2184
rect 7332 -2242 7384 -2236
rect 7943 -2239 7952 -2235
rect 8012 -2239 8021 -2179
rect 8114 -2353 8166 -2128
rect 9104 -2076 9156 -2070
rect 9104 -2134 9156 -2128
rect 10114 -2072 10166 -2066
rect 11008 -2076 11055 -1805
rect 11258 -1990 11298 -1800
rect 11701 -1957 11745 -1650
rect 12142 -1743 12187 -1195
rect 12275 -1226 12327 -1220
rect 12712 -1262 12750 -966
rect 13143 -1140 13193 -799
rect 13702 -986 13708 -934
rect 13760 -986 13766 -934
rect 13142 -1146 13194 -1140
rect 13142 -1204 13194 -1198
rect 12275 -1284 12327 -1278
rect 12282 -1604 12319 -1284
rect 12686 -1314 12692 -1262
rect 12770 -1314 12776 -1262
rect 12282 -1641 12750 -1604
rect 12142 -1788 12310 -1743
rect 11252 -1996 11304 -1990
rect 11678 -2009 11684 -1957
rect 11762 -2009 11768 -1957
rect 12265 -1981 12310 -1788
rect 12713 -1955 12750 -1641
rect 13143 -1739 13193 -1204
rect 13274 -1222 13326 -1216
rect 13714 -1230 13754 -986
rect 14143 -1131 14192 -650
rect 14879 -660 14888 -604
rect 14944 -660 14953 -604
rect 14886 -1034 14946 -660
rect 14142 -1137 14194 -1131
rect 14895 -1175 14938 -1034
rect 15173 -1130 15223 -481
rect 15587 -486 15639 -480
rect 16601 -544 16639 528
rect 16724 515 16767 718
rect 17584 520 17590 572
rect 17668 520 17674 572
rect 16720 509 16772 515
rect 16720 451 16772 457
rect 16588 -596 16594 -544
rect 16646 -596 16652 -544
rect 17609 -692 17649 520
rect 17734 509 17777 718
rect 17730 503 17782 509
rect 17730 445 17782 451
rect 17603 -698 17655 -692
rect 17603 -756 17655 -750
rect 18691 -861 18741 861
rect 15313 -911 18741 -861
rect 15172 -1136 15224 -1130
rect 14142 -1195 14194 -1189
rect 13274 -1280 13326 -1274
rect 13708 -1236 13760 -1230
rect 13280 -1604 13320 -1280
rect 13708 -1294 13760 -1288
rect 13280 -1644 13759 -1604
rect 13143 -1789 13319 -1739
rect 12262 -1987 12314 -1981
rect 12686 -2007 12692 -1955
rect 12770 -2007 12776 -1955
rect 13272 -1988 13316 -1789
rect 13719 -1961 13759 -1644
rect 14143 -1737 14192 -1195
rect 14289 -1228 14341 -1222
rect 14289 -1286 14341 -1280
rect 14293 -1609 14336 -1286
rect 14293 -1652 14769 -1609
rect 14143 -1786 14330 -1737
rect 13268 -1994 13320 -1988
rect 12262 -2045 12314 -2039
rect 11252 -2054 11304 -2048
rect 13694 -2013 13700 -1961
rect 13778 -2013 13784 -1961
rect 14281 -1981 14330 -1786
rect 14726 -1967 14769 -1652
rect 14280 -1987 14332 -1981
rect 14702 -2019 14708 -1967
rect 14786 -2019 14792 -1967
rect 14280 -2045 14332 -2039
rect 13268 -2052 13320 -2046
rect 11126 -2076 11132 -2073
rect 11008 -2123 11132 -2076
rect 10114 -2130 10166 -2124
rect 11126 -2125 11132 -2123
rect 11184 -2125 11190 -2073
rect 12140 -2074 12192 -2068
rect 12140 -2132 12192 -2126
rect 8114 -2411 8166 -2405
rect 9109 -2438 9151 -2134
rect 9576 -2180 9632 -2171
rect 12142 -2184 12189 -2132
rect 13138 -2134 13144 -2082
rect 13196 -2089 13202 -2082
rect 13196 -2134 13264 -2089
rect 14145 -2121 14151 -2069
rect 14203 -2075 14209 -2069
rect 14896 -2075 14937 -1175
rect 15172 -1194 15224 -1188
rect 15155 -1598 15215 -1589
rect 15153 -1654 15155 -1602
rect 15215 -1654 15217 -1602
rect 15155 -1667 15215 -1658
rect 14203 -2116 14937 -2075
rect 14203 -2121 14209 -2116
rect 13198 -2160 13264 -2134
rect 9632 -2231 12189 -2184
rect 9576 -2245 9632 -2236
rect 13226 -2296 13264 -2160
rect 13127 -2352 13136 -2296
rect 13192 -2351 13273 -2296
rect 13192 -2352 13201 -2351
rect -17 -2511 7278 -2461
rect 9102 -2488 9158 -2438
rect 15316 -2483 15361 -911
rect 15307 -2535 15313 -2483
rect 15365 -2535 15371 -2483
rect 9102 -2553 9158 -2544
<< via2 >>
rect 323 40 383 100
rect 7144 -34 7200 22
rect 9158 -474 9218 -414
rect 3310 -894 3370 -834
rect 6918 -954 6978 -894
rect 3356 -1573 3416 -1513
rect 10368 -144 10428 -84
rect 15008 -30 15064 26
rect 3922 -1540 3978 -1484
rect 5608 -1554 5664 -1502
rect 5608 -1558 5664 -1554
rect 5606 -1764 5666 -1704
rect 5902 -1767 5962 -1707
rect 6426 -1862 6430 -1812
rect 6430 -1862 6482 -1812
rect 6426 -1868 6482 -1862
rect 12136 -952 12192 -896
rect 11128 -1128 11184 -1072
rect 6612 -2409 6672 -2349
rect 6904 -2407 6960 -2351
rect 10030 -1970 10086 -1914
rect 7952 -2239 8012 -2179
rect 14888 -660 14944 -604
rect 9576 -2236 9632 -2180
rect 15155 -1602 15215 -1598
rect 15155 -1654 15159 -1602
rect 15159 -1654 15211 -1602
rect 15211 -1654 15215 -1602
rect 15155 -1658 15215 -1654
rect 13136 -2352 13192 -2296
rect 9102 -2544 9158 -2488
<< metal3 >>
rect 318 100 388 105
rect -26 40 323 100
rect 383 40 388 100
rect -26 -2486 34 40
rect 318 35 388 40
rect 15003 28 15069 31
rect 15153 30 15217 36
rect 7139 22 7205 27
rect 7139 -34 7144 22
rect 7200 -34 7205 22
rect 7139 -38 7205 -34
rect 15003 26 15153 28
rect 15003 -30 15008 26
rect 15064 -30 15153 26
rect 15003 -32 15153 -30
rect 15003 -35 15069 -32
rect 7139 -39 7208 -38
rect 7142 -84 7208 -39
rect 15153 -40 15217 -34
rect 10363 -84 10433 -79
rect 7142 -144 10368 -84
rect 10428 -144 10433 -84
rect 10363 -149 10433 -144
rect 9153 -414 9223 -409
rect 9153 -474 9158 -414
rect 9218 -474 14946 -414
rect 9153 -479 9223 -474
rect 14886 -599 14946 -474
rect 14883 -604 14949 -599
rect 14883 -660 14888 -604
rect 14944 -660 14949 -604
rect 14883 -665 14949 -660
rect 3305 -834 3375 -829
rect 3305 -894 3310 -834
rect 3370 -894 6594 -834
rect 3305 -899 3375 -894
rect 3917 -1484 3983 -1479
rect 6534 -1484 6594 -894
rect 6913 -894 6983 -889
rect 12131 -894 12197 -891
rect 6913 -954 6918 -894
rect 6978 -896 12197 -894
rect 6978 -952 12136 -896
rect 12192 -952 12197 -896
rect 6978 -954 12197 -952
rect 6913 -959 6983 -954
rect 12131 -957 12197 -954
rect 11123 -1070 11189 -1067
rect 6762 -1072 11189 -1070
rect 6762 -1128 11128 -1072
rect 11184 -1128 11189 -1072
rect 6762 -1130 11189 -1128
rect 3351 -1513 3421 -1508
rect 3917 -1513 3922 -1484
rect 3351 -1573 3356 -1513
rect 3416 -1540 3922 -1513
rect 3978 -1540 3983 -1484
rect 3416 -1545 3983 -1540
rect 5603 -1502 5669 -1497
rect 3416 -1573 3980 -1545
rect 5603 -1558 5608 -1502
rect 5664 -1558 5669 -1502
rect 6526 -1548 6532 -1484
rect 6596 -1548 6602 -1484
rect 5603 -1563 5669 -1558
rect 3351 -1578 3421 -1573
rect 5606 -1699 5666 -1563
rect 6762 -1618 6822 -1130
rect 11123 -1133 11189 -1130
rect 15153 -1408 15217 -1402
rect 15153 -1478 15217 -1472
rect 15155 -1593 15215 -1478
rect 6424 -1678 6822 -1618
rect 15150 -1598 15220 -1593
rect 15150 -1658 15155 -1598
rect 15215 -1658 15220 -1598
rect 15150 -1663 15220 -1658
rect 5601 -1704 5671 -1699
rect 5601 -1764 5606 -1704
rect 5666 -1764 5671 -1704
rect 5601 -1769 5671 -1764
rect 5897 -1707 5967 -1702
rect 5897 -1767 5902 -1707
rect 5962 -1767 5967 -1707
rect 5897 -1772 5967 -1767
rect 5902 -2200 5962 -1772
rect 6424 -1807 6484 -1678
rect 6421 -1812 6487 -1807
rect 6421 -1868 6426 -1812
rect 6482 -1868 6487 -1812
rect 6421 -1873 6487 -1868
rect 10025 -1912 10091 -1909
rect 9896 -1914 10091 -1912
rect 9896 -1970 10030 -1914
rect 10086 -1970 10091 -1914
rect 9896 -1972 10091 -1970
rect 9896 -2070 9956 -1972
rect 10025 -1975 10091 -1972
rect 9894 -2076 9958 -2070
rect 9894 -2146 9958 -2140
rect 7947 -2179 8017 -2174
rect 9571 -2178 9637 -2175
rect 9210 -2179 9637 -2178
rect 5900 -2206 5964 -2200
rect 7947 -2239 7952 -2179
rect 8012 -2180 9637 -2179
rect 8012 -2236 9576 -2180
rect 9632 -2236 9637 -2180
rect 8012 -2239 9637 -2236
rect 7947 -2244 8017 -2239
rect 9571 -2241 9637 -2239
rect 5900 -2276 5964 -2270
rect 13131 -2296 13197 -2291
rect 6607 -2349 6677 -2344
rect 6899 -2349 6965 -2346
rect 6607 -2409 6612 -2349
rect 6672 -2351 6965 -2349
rect 6672 -2407 6904 -2351
rect 6960 -2407 6965 -2351
rect 13131 -2352 13136 -2296
rect 13192 -2352 13197 -2296
rect 13131 -2357 13197 -2352
rect 6672 -2409 6965 -2407
rect 6607 -2414 6677 -2409
rect 6899 -2412 6965 -2409
rect 13134 -2436 13194 -2357
rect 13132 -2442 13196 -2436
rect 9097 -2486 9163 -2483
rect -26 -2488 9163 -2486
rect -26 -2544 9102 -2488
rect 9158 -2544 9163 -2488
rect 13132 -2512 13196 -2506
rect -26 -2546 9163 -2544
rect 9097 -2549 9163 -2546
<< via3 >>
rect 15153 -34 15217 30
rect 6532 -1548 6596 -1484
rect 15153 -1472 15217 -1408
rect 9894 -2140 9958 -2076
rect 5900 -2270 5964 -2206
rect 13132 -2506 13196 -2442
<< metal4 >>
rect 15152 30 15218 31
rect 15152 -34 15153 30
rect 15217 -34 15218 30
rect 15152 -35 15218 -34
rect 15155 -1407 15215 -35
rect 15152 -1408 15218 -1407
rect 15152 -1472 15153 -1408
rect 15217 -1472 15218 -1408
rect 15152 -1473 15218 -1472
rect 6531 -1484 6597 -1483
rect 6531 -1548 6532 -1484
rect 6596 -1548 6597 -1484
rect 6531 -1549 6597 -1548
rect 6534 -2078 6594 -1549
rect 9893 -2076 9959 -2075
rect 9893 -2078 9894 -2076
rect 6534 -2138 9894 -2078
rect 9893 -2140 9894 -2138
rect 9958 -2140 9959 -2076
rect 9893 -2141 9959 -2140
rect 5899 -2206 5965 -2205
rect 5899 -2270 5900 -2206
rect 5964 -2270 5965 -2206
rect 5899 -2271 5965 -2270
rect 5902 -2444 5962 -2271
rect 13131 -2442 13197 -2441
rect 13131 -2444 13132 -2442
rect 5902 -2504 13132 -2444
rect 13131 -2506 13132 -2504
rect 13196 -2506 13197 -2442
rect 13131 -2507 13197 -2506
use DFF  DFF_0
timestamp 1681866284
transform 1 0 234 0 1 46
box -268 0 3242 976
use DFF  DFF_1
timestamp 1681866284
transform 1 0 234 0 -1 142
box -268 0 3242 976
use DFF  DFF_2
timestamp 1681866284
transform 1 0 234 0 -1 -1586
box -268 0 3242 976
use DFF  DFF_3
timestamp 1681866284
transform 1 0 234 0 1 -1682
box -268 0 3242 976
use DFF  DFF_4
timestamp 1681866284
transform 1 0 3686 0 1 -1682
box -268 0 3242 976
use DFF  DFF_5
timestamp 1681866284
transform 1 0 3686 0 -1 -1586
box -268 0 3242 976
use DFF  DFF_6
timestamp 1681866284
transform 1 0 3686 0 -1 142
box -268 0 3242 976
use DFF  DFF_7
timestamp 1681866284
transform 1 0 3686 0 1 46
box -268 0 3242 976
use DFF  DFF_8
timestamp 1681866284
transform 1 0 7138 0 1 46
box -268 0 3242 976
use multiplexor  multiplexor_0
timestamp 1681434240
transform 1 0 7138 0 1 -1682
box -268 0 8162 976
use multiplexor  multiplexor_1
timestamp 1681434240
transform 1 0 7138 0 -1 -1586
box -268 0 8162 976
use multiplexor  multiplexor_2
timestamp 1681434240
transform 1 0 10590 0 1 46
box -268 0 8162 976
<< labels >>
flabel locali s 48 444 114 510 0 FreeSerif 800 0 0 0 CLK
port 0 nsew
flabel locali s 10404 444 10470 510 0 FreeSerif 800 0 0 0 A
port 10 nsew
flabel locali s 18166 374 18232 676 0 FreeSerif 800 0 0 0 Y7
port 22 nsew
flabel locali s 17158 374 17224 676 0 FreeSerif 800 0 0 0 Y6
port 21 nsew
flabel locali s 16150 374 16216 676 0 FreeSerif 800 0 0 0 Y5
port 20 nsew
flabel locali s 15142 374 15208 676 0 FreeSerif 800 0 0 0 Y4
port 19 nsew
flabel locali s 14134 374 14200 676 0 FreeSerif 800 0 0 0 Y3
port 18 nsew
flabel locali s 13126 374 13192 676 0 FreeSerif 800 0 0 0 Y2
port 17 nsew
flabel locali s 12118 374 12184 676 0 FreeSerif 800 0 0 0 Y1
port 16 nsew
flabel locali s 11110 374 11176 676 0 FreeSerif 800 0 0 0 Y0
port 15 nsew
flabel locali s 6952 -1284 7018 -1218 0 FreeSerif 800 0 0 0 B
port 11 nsew
flabel locali s -30 -2546 15296 -2450 0 FreeSerif 1600 0 0 0 VDD!
flabel locali s -30 -1682 15296 -1586 0 FreeSerif 1600 0 0 0 GND!
<< end >>
