magic
tech sky130A
timestamp 1677800174
<< nwell >>
rect -42 135 283 426
<< nmos >>
rect 32 3 47 53
rect 68 3 83 53
rect 122 3 137 53
rect 158 3 173 53
<< pmos >>
rect 32 219 47 319
rect 86 219 101 319
rect 140 219 155 319
rect 194 219 209 319
<< ndiff >>
rect -7 45 32 53
rect -7 11 4 45
rect 21 11 32 45
rect -7 3 32 11
rect 47 3 68 53
rect 83 45 122 53
rect 83 11 94 45
rect 111 11 122 45
rect 83 3 122 11
rect 137 3 158 53
rect 173 45 212 53
rect 173 11 184 45
rect 201 11 212 45
rect 173 3 212 11
<< pdiff >>
rect -4 311 32 319
rect -4 227 4 311
rect 21 227 32 311
rect -4 219 32 227
rect 47 311 86 319
rect 47 227 58 311
rect 75 227 86 311
rect 47 219 86 227
rect 101 311 140 319
rect 101 227 112 311
rect 129 227 140 311
rect 101 219 140 227
rect 155 311 194 319
rect 155 227 166 311
rect 183 227 194 311
rect 155 219 194 227
rect 209 311 248 319
rect 209 227 220 311
rect 237 227 248 311
rect 209 219 248 227
<< ndiffc >>
rect 4 11 21 45
rect 94 11 111 45
rect 184 11 201 45
<< pdiffc >>
rect 4 227 21 311
rect 58 227 75 311
rect 112 227 129 311
rect 166 227 183 311
rect 220 227 237 311
<< psubdiff >>
rect -4 -52 8 -24
rect 111 -52 123 -24
<< nsubdiff >>
rect 3 380 15 408
rect 118 380 130 408
<< psubdiffcont >>
rect 8 -52 111 -24
<< nsubdiffcont >>
rect 15 380 118 408
<< poly >>
rect 32 319 47 332
rect 86 319 101 332
rect 140 319 155 332
rect 194 319 209 332
rect 32 210 47 219
rect 10 195 47 210
rect 10 161 25 195
rect -23 153 25 161
rect 86 154 101 219
rect -23 136 -15 153
rect 2 136 25 153
rect -23 128 25 136
rect 10 79 25 128
rect 53 146 101 154
rect 53 129 61 146
rect 78 129 101 146
rect 53 121 101 129
rect 86 79 101 121
rect 140 133 155 219
rect 194 190 209 219
rect 194 175 224 190
rect 140 125 188 133
rect 140 115 163 125
rect 10 64 47 79
rect 32 53 47 64
rect 68 64 101 79
rect 122 108 163 115
rect 180 108 188 125
rect 122 100 188 108
rect 209 106 224 175
rect 68 53 83 64
rect 122 53 137 100
rect 209 98 257 106
rect 209 81 232 98
rect 249 81 257 98
rect 209 79 257 81
rect 158 73 257 79
rect 158 64 224 73
rect 158 53 173 64
rect 32 -10 47 3
rect 68 -10 83 3
rect 122 -10 137 3
rect 158 -10 173 3
<< polycont >>
rect -15 136 2 153
rect 61 129 78 146
rect 163 108 180 125
rect 232 81 249 98
<< locali >>
rect -40 408 281 418
rect -40 380 15 408
rect 118 380 281 408
rect -40 370 281 380
rect -4 311 29 319
rect -4 227 4 311
rect 21 227 29 311
rect -4 201 29 227
rect 50 311 83 370
rect 50 227 58 311
rect 75 227 83 311
rect 50 219 83 227
rect 104 336 245 353
rect 104 311 137 336
rect 104 227 112 311
rect 129 227 137 311
rect 104 201 137 227
rect -4 188 137 201
rect 158 311 191 319
rect 158 227 166 311
rect 183 227 191 311
rect -4 184 121 188
rect -4 179 105 184
rect 158 171 191 227
rect 212 311 245 336
rect 212 227 220 311
rect 237 227 245 311
rect 212 219 245 227
rect 136 167 191 171
rect 120 162 191 167
rect -23 153 10 161
rect 111 154 191 162
rect -23 136 -15 153
rect 2 136 10 153
rect -23 128 10 136
rect 53 146 86 154
rect 53 129 61 146
rect 78 129 86 146
rect 53 121 86 129
rect 111 150 155 154
rect 111 104 137 150
rect 86 83 137 104
rect 155 125 188 133
rect 155 108 163 125
rect 180 108 188 125
rect 155 100 188 108
rect 224 98 257 106
rect -4 45 29 53
rect -4 11 4 45
rect 21 11 29 45
rect -4 -14 29 11
rect 86 45 119 83
rect 224 81 232 98
rect 249 81 257 98
rect 224 73 257 81
rect 86 11 94 45
rect 111 11 119 45
rect 86 3 119 11
rect 176 45 209 53
rect 176 11 184 45
rect 201 11 209 45
rect 176 -14 209 11
rect -40 -24 281 -14
rect -40 -52 8 -24
rect 111 -52 281 -24
rect -40 -62 281 -52
<< labels >>
flabel locali -40 370 281 418 0 FreeSerif 80 0 0 0 VDD!
port 0 nsew
flabel locali -40 -62 281 -14 0 FreeSerif 80 0 0 0 GND!
port 1 nsew
flabel locali 53 121 86 154 0 FreeSerif 80 0 0 0 A
port 11 nsew
flabel locali -23 128 10 161 0 FreeSerif 80 0 0 0 B
port 12 nsew
flabel locali 158 154 191 219 0 FreeSerif 80 0 0 0 Y
port 4 nsew
flabel locali 155 100 188 133 0 FreeSerif 80 0 0 0 NOT_B
port 14 nsew
flabel locali 224 73 257 106 0 FreeSerif 80 0 0 0 NOT_A
port 13 nsew
<< end >>
