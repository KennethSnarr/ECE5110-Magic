magic
tech sky130A
magscale 1 2
timestamp 1681869295
<< locali >>
rect 4 1728 13866 1824
rect 3004 1591 3070 1594
rect 3004 1430 3070 1551
rect 3340 1430 3406 1561
rect 6456 1593 6522 1594
rect 6456 1430 6522 1559
rect 6792 1593 6858 1594
rect 6792 1430 6858 1559
rect 9908 1593 9974 1594
rect 9908 1430 9974 1551
rect 10244 1430 10310 1561
rect 13360 1430 13426 1594
rect 13696 1430 13762 1594
rect -3448 864 13866 960
rect -3102 528 -3036 594
rect -3376 386 -3304 476
rect -448 274 -382 394
rect -448 230 -382 231
rect -112 263 -46 394
rect 76 386 148 476
rect 3004 297 3070 394
rect 3004 231 3029 297
rect 3004 230 3070 231
rect 3340 276 3406 394
rect 3528 386 3600 476
rect 3340 230 3406 235
rect 6456 276 6522 394
rect 6456 230 6522 233
rect 6792 275 6858 394
rect 6792 230 6858 233
rect 9908 272 9974 394
rect 9908 230 9974 231
rect 10244 276 10310 394
rect 13360 265 13426 394
rect 13360 230 13426 231
rect 13696 271 13762 394
rect 13696 230 13762 231
rect -3448 0 13866 96
<< viali >>
rect 3004 1551 3070 1591
rect 3340 1561 3406 1595
rect 6456 1559 6522 1593
rect 6792 1559 6858 1593
rect 9908 1551 9974 1593
rect 10244 1561 10310 1595
rect -448 231 -382 274
rect -112 229 -46 263
rect 3029 231 3070 297
rect 3340 235 3406 276
rect 6456 233 6522 276
rect 6792 233 6858 275
rect 9908 231 9974 272
rect 10244 229 10310 276
rect 13360 231 13426 265
rect 13696 231 13762 271
<< metal1 >>
rect 3017 1668 3586 1708
rect 3017 1597 3057 1668
rect 3334 1604 3412 1610
rect 2992 1591 3082 1597
rect 2992 1551 3004 1591
rect 3070 1551 3082 1591
rect 3328 1555 3334 1601
rect 2992 1545 3082 1551
rect 3412 1555 3418 1601
rect 3334 1546 3412 1552
rect 85 880 116 1423
rect 3546 1374 3586 1668
rect 6472 1659 7033 1693
rect 6472 1599 6506 1659
rect 6786 1602 6864 1608
rect 6444 1593 6534 1599
rect 6444 1559 6456 1593
rect 6522 1559 6534 1593
rect 6444 1553 6534 1559
rect 6780 1553 6786 1599
rect 6864 1553 6870 1599
rect 6786 1544 6864 1550
rect 6999 1381 7033 1659
rect 9920 1659 10489 1701
rect 9920 1599 9962 1659
rect 10238 1604 10316 1610
rect 9896 1593 9986 1599
rect 9896 1551 9908 1593
rect 9974 1551 9986 1593
rect 10232 1555 10238 1601
rect 9896 1545 9986 1551
rect 10316 1555 10322 1601
rect 10238 1546 10316 1552
rect 10447 1375 10489 1659
rect 363 947 393 1287
rect 3347 1007 3399 1013
rect 3346 955 3347 956
rect 3346 949 3399 955
rect 3813 967 3844 1271
rect 6800 977 6852 983
rect 3346 947 3388 949
rect 363 917 3388 947
rect 3813 936 6800 967
rect 7261 957 7292 1285
rect 10246 957 10252 967
rect 7261 926 10252 957
rect 6800 919 6852 925
rect 10246 915 10252 926
rect 10304 915 10310 967
rect 13368 890 13420 896
rect 85 849 13368 880
rect 13368 832 13420 838
rect -3096 540 -3090 592
rect -3038 540 -3032 592
rect 344 540 350 592
rect 402 540 408 592
rect 3800 536 3806 588
rect 3858 536 3864 588
rect 7246 522 7252 574
rect 7304 522 7310 574
rect 10704 534 10710 586
rect 10762 534 10768 586
rect 92 410 98 462
rect 150 410 156 462
rect 3542 414 3548 466
rect 3600 414 3606 466
rect 6986 412 6992 464
rect 7044 412 7050 464
rect 10440 408 10446 460
rect 10498 408 10504 460
rect 3023 303 3076 309
rect -454 280 -376 283
rect -460 277 -370 280
rect -460 225 -454 277
rect -376 225 -370 277
rect -124 263 -34 269
rect -124 229 -112 263
rect -46 229 -34 263
rect -454 219 -376 225
rect -124 223 -34 229
rect 3018 225 3024 303
rect 3076 225 3082 303
rect 6450 282 6528 285
rect 3328 276 3418 282
rect 3328 235 3340 276
rect 3406 235 3418 276
rect 3328 229 3418 235
rect 6444 279 6534 282
rect -96 100 -62 223
rect 3023 219 3076 225
rect -111 48 -105 100
rect -53 48 -47 100
rect 343 43 349 95
rect 401 89 407 95
rect 3353 89 3394 229
rect 6444 227 6450 279
rect 6528 227 6534 279
rect 6780 275 6870 281
rect 9902 278 9980 283
rect 6780 233 6792 275
rect 6858 233 6870 275
rect 6780 227 6870 233
rect 9896 277 9986 278
rect 6450 221 6528 227
rect 401 48 3394 89
rect 3806 88 3858 94
rect 401 43 407 48
rect 6804 83 6846 227
rect 9896 225 9902 277
rect 9980 225 9986 277
rect 10232 276 10322 282
rect 10232 229 10244 276
rect 10310 229 10322 276
rect 13354 274 13432 280
rect 9902 219 9980 225
rect 10232 223 10322 229
rect 13348 225 13354 271
rect 13684 271 13774 277
rect 3858 41 6846 83
rect 7251 89 7303 95
rect 3806 30 3858 36
rect 10254 83 10301 223
rect 13432 225 13438 271
rect 13684 231 13696 271
rect 13762 231 13774 271
rect 13684 225 13774 231
rect 13354 216 13432 222
rect 7303 42 10301 83
rect 10254 39 10301 42
rect 10710 84 10762 90
rect 7251 31 7303 37
rect 13709 76 13749 225
rect 10762 40 13749 76
rect 13709 38 13749 40
rect 10710 26 10762 32
<< via1 >>
rect 3334 1595 3412 1604
rect 3334 1561 3340 1595
rect 3340 1561 3406 1595
rect 3406 1561 3412 1595
rect 3334 1552 3412 1561
rect 6786 1593 6864 1602
rect 6786 1559 6792 1593
rect 6792 1559 6858 1593
rect 6858 1559 6864 1593
rect 6786 1550 6864 1559
rect 10238 1595 10316 1604
rect 10238 1561 10244 1595
rect 10244 1561 10310 1595
rect 10310 1561 10316 1595
rect 10238 1552 10316 1561
rect 3347 955 3399 1007
rect 6800 925 6852 977
rect 10252 915 10304 967
rect 13368 838 13420 890
rect -3090 540 -3038 592
rect 350 540 402 592
rect 3806 536 3858 588
rect 7252 522 7304 574
rect 10710 534 10762 586
rect 98 410 150 462
rect 3548 414 3600 466
rect 6992 412 7044 464
rect 10446 408 10498 460
rect -454 274 -376 277
rect -454 231 -448 274
rect -448 231 -382 274
rect -382 231 -376 274
rect -454 225 -376 231
rect 3024 297 3076 303
rect 3024 231 3029 297
rect 3029 231 3070 297
rect 3070 231 3076 297
rect 3024 225 3076 231
rect -105 48 -53 100
rect 349 43 401 95
rect 6450 276 6528 279
rect 6450 233 6456 276
rect 6456 233 6522 276
rect 6522 233 6528 276
rect 6450 227 6528 233
rect 3806 36 3858 88
rect 9902 272 9980 277
rect 9902 231 9908 272
rect 9908 231 9974 272
rect 9974 231 9980 272
rect 9902 225 9980 231
rect 13354 265 13432 274
rect 13354 231 13360 265
rect 13360 231 13426 265
rect 13426 231 13432 265
rect 7251 37 7303 89
rect 13354 222 13432 231
rect 10710 32 10762 84
<< metal2 >>
rect 3328 1552 3334 1604
rect 3412 1552 3418 1604
rect 3358 1007 3388 1552
rect 6780 1550 6786 1602
rect 6864 1550 6870 1602
rect 10232 1552 10238 1604
rect 10316 1552 10322 1604
rect 3341 955 3347 1007
rect 3399 955 3405 1007
rect 6810 977 6841 1550
rect 6794 925 6800 977
rect 6852 925 6858 977
rect 10262 973 10293 1552
rect 10252 967 10304 973
rect 10252 909 10304 915
rect 13362 838 13368 890
rect 13420 838 13426 890
rect -3090 592 -3038 598
rect -3090 534 -3038 540
rect 350 592 402 598
rect 350 534 402 540
rect 3806 588 3858 594
rect 10710 586 10762 592
rect -3081 91 -3047 534
rect 98 462 150 468
rect 98 404 150 410
rect -460 225 -454 277
rect -376 274 -370 277
rect 101 274 146 404
rect -376 229 146 274
rect -376 225 -370 229
rect -105 100 -53 106
rect 355 101 396 534
rect 3806 530 3858 536
rect 7252 574 7304 580
rect 3548 466 3600 472
rect 3548 408 3600 414
rect 3024 303 3076 309
rect 3553 285 3594 408
rect 3076 244 3594 285
rect 3024 219 3076 225
rect -3081 57 -105 91
rect -105 42 -53 48
rect 349 95 401 101
rect 3811 88 3853 530
rect 10710 528 10762 534
rect 7252 516 7304 522
rect 6992 464 7044 470
rect 6992 406 7044 412
rect 6444 227 6450 279
rect 6528 275 6534 279
rect 6996 275 7039 406
rect 6528 232 7039 275
rect 6528 227 6534 232
rect 7257 89 7298 516
rect 10446 460 10498 466
rect 10446 402 10498 408
rect 9896 225 9902 277
rect 9980 272 9986 277
rect 10451 272 10492 402
rect 9980 231 10492 272
rect 9980 225 9986 231
rect 349 37 401 43
rect 3800 36 3806 88
rect 3858 36 3864 88
rect 7245 37 7251 89
rect 7303 37 7309 89
rect 10718 84 10754 528
rect 13378 274 13409 838
rect 13348 222 13354 274
rect 13432 222 13438 274
rect 10704 32 10710 84
rect 10762 32 10768 84
use DFF  DFF_0
timestamp 1681866284
transform 1 0 268 0 1 0
box -268 0 3242 976
use DFF  DFF_1
timestamp 1681866284
transform 1 0 3720 0 1 0
box -268 0 3242 976
use DFF  DFF_2
timestamp 1681866284
transform 1 0 7172 0 1 0
box -268 0 3242 976
use DFF  DFF_3
timestamp 1681866284
transform 1 0 10624 0 1 0
box -268 0 3242 976
use DFF  DFF_4
timestamp 1681866284
transform 1 0 10624 0 -1 1824
box -268 0 3242 976
use DFF  DFF_5
timestamp 1681866284
transform 1 0 7172 0 -1 1824
box -268 0 3242 976
use DFF  DFF_6
timestamp 1681866284
transform 1 0 3720 0 -1 1824
box -268 0 3242 976
use DFF  DFF_7
timestamp 1681866284
transform 1 0 268 0 -1 1824
box -268 0 3242 976
use DFF  DFF_8
timestamp 1681866284
transform 1 0 -3184 0 1 0
box -268 0 3242 976
<< labels >>
flabel locali s -3376 386 -3304 476 0 FreeSerif 560 0 0 0 CLK
<< end >>
