magic
tech sky130A
magscale 1 2
timestamp 1680050683
<< poly >>
rect 3756 104 3786 106
<< locali >>
rect 4 864 4184 960
rect 1680 612 1746 630
rect 976 514 1042 562
rect 82 396 148 464
rect 390 398 456 466
rect 976 461 982 514
rect 1035 461 1042 514
rect 976 432 1042 461
rect 1680 560 1686 612
rect 1738 560 1746 612
rect 1680 230 1746 560
rect 2126 398 2192 464
rect 2712 432 2778 562
rect 3416 327 3482 630
rect 3587 398 3648 464
rect 3684 458 3750 542
rect 3684 404 3689 458
rect 3743 404 3750 458
rect 3416 273 3421 327
rect 3475 273 3482 327
rect 3416 230 3482 273
rect 3684 230 3750 404
rect 3786 333 3852 382
rect 4046 230 4112 630
rect 4 0 4184 96
<< viali >>
rect 982 461 1035 514
rect 1686 560 1738 612
rect 1818 398 1884 464
rect 3521 398 3587 464
rect 3689 404 3743 458
rect 3421 273 3475 327
rect 3944 398 4010 464
rect 3786 267 3852 333
<< metal1 >>
rect 1680 700 3586 764
rect 1680 612 1744 700
rect 1680 560 1686 612
rect 1738 560 1744 612
rect 1680 548 1744 560
rect 976 520 1041 526
rect 3522 476 3586 700
rect 976 449 1041 455
rect 1806 392 1812 470
rect 1877 464 1896 470
rect 1884 398 1896 464
rect 1877 392 1896 398
rect 3515 464 3593 476
rect 3938 464 4016 476
rect 3515 398 3521 464
rect 3587 398 3593 464
rect 3677 458 3944 464
rect 3677 404 3689 458
rect 3743 404 3944 458
rect 3677 398 3944 404
rect 4010 398 4016 464
rect 3515 386 3593 398
rect 3938 386 4016 398
rect 3774 333 3864 339
rect 3409 327 3786 333
rect 3409 273 3421 327
rect 3475 273 3786 327
rect 3409 267 3786 273
rect 3852 267 3864 333
rect 3774 261 3864 267
<< via1 >>
rect 976 514 1041 520
rect 976 461 982 514
rect 982 461 1035 514
rect 1035 461 1041 514
rect 976 455 1041 461
rect 1812 464 1877 470
rect 1812 398 1818 464
rect 1818 398 1877 464
rect 1812 392 1877 398
<< metal2 >>
rect 970 455 976 520
rect 1041 464 1175 520
rect 1812 470 1877 476
rect 1041 455 1812 464
rect 1110 399 1812 455
rect 1812 386 1877 392
use half_adder  half_adder_0
timestamp 1679945325
transform 1 0 576 0 1 0
box -576 0 1246 976
use half_adder  half_adder_1
timestamp 1679945325
transform 1 0 2312 0 1 0
box -576 0 1246 976
use inv  inv_0
timestamp 1679616770
transform 1 0 3946 0 1 124
box -84 -124 242 852
use nor2  nor2_0
timestamp 1676660012
transform 1 0 3584 0 1 124
box -84 -124 350 852
<< labels >>
flabel locali 82 396 148 464 0 FreeSerif 240 0 0 0 A
port 1 nsew
flabel locali 390 398 456 466 0 FreeSerif 240 0 0 0 B
port 2 nsew
flabel locali s 4046 230 4112 630 0 FreeSerif 240 0 0 0 C_out
port 3 nsew
flabel locali s 2712 432 2778 562 0 FreeSerif 240 0 0 0 S
port 0 nsew
<< end >>
