magic
tech sky130A
timestamp 1679945325
<< poly >>
rect 422 265 455 273
rect 422 248 430 265
rect 447 248 455 265
rect 422 240 455 248
rect -247 224 -214 232
rect -247 207 -239 224
rect -222 207 -214 224
rect -247 199 -214 207
rect -93 224 -60 232
rect -93 207 -85 224
rect -68 207 -60 224
rect 320 224 353 232
rect -93 199 -60 207
rect 19 215 52 223
rect 19 198 27 215
rect 44 198 52 215
rect 19 190 52 198
rect 95 208 128 216
rect 95 191 103 208
rect 120 191 128 208
rect 320 207 328 224
rect 345 207 353 224
rect 320 199 353 207
rect 501 224 534 232
rect 501 207 509 224
rect 526 207 534 224
rect 501 199 534 207
rect 95 183 128 191
rect 197 187 230 195
rect 197 170 205 187
rect 222 170 230 187
rect 197 162 230 170
rect 266 160 299 168
rect 266 143 274 160
rect 291 143 299 160
rect 266 135 299 143
<< polycont >>
rect 430 248 447 265
rect -239 207 -222 224
rect -85 207 -68 224
rect 27 198 44 215
rect 103 191 120 208
rect 328 207 345 224
rect 509 207 526 224
rect 205 170 222 187
rect 274 143 291 160
<< locali >>
rect -286 432 621 480
rect -247 224 -214 232
rect -247 207 -239 224
rect -222 207 -214 224
rect -247 199 -214 207
rect -196 109 -163 315
rect -93 224 -60 232
rect -93 207 -85 224
rect -68 207 -60 224
rect -93 199 -60 207
rect -42 138 -9 315
rect 371 306 404 315
rect 371 289 378 306
rect 396 289 404 306
rect 19 215 52 223
rect 200 216 233 281
rect 320 224 353 232
rect 19 198 27 215
rect 44 198 52 215
rect 19 190 52 198
rect 95 208 128 216
rect 95 191 103 208
rect 120 191 128 208
rect 320 207 328 224
rect 345 207 353 224
rect 320 199 353 207
rect 95 183 128 191
rect 197 187 230 195
rect 197 170 205 187
rect 222 170 230 187
rect 197 162 230 170
rect -42 121 -35 138
rect -18 121 -9 138
rect 266 160 299 168
rect 371 164 404 289
rect 422 265 455 273
rect 422 248 430 265
rect 447 248 455 265
rect 422 240 455 248
rect 501 224 534 232
rect 501 207 509 224
rect 526 207 534 224
rect 501 199 534 207
rect 266 143 274 160
rect 291 143 299 160
rect 266 135 299 143
rect -42 115 -9 121
rect 552 115 585 315
rect -196 87 -191 109
rect -169 87 -163 109
rect -196 82 -163 87
rect -286 0 621 48
<< viali >>
rect -239 207 -222 224
rect -85 207 -68 224
rect 378 289 396 306
rect 27 198 44 215
rect 103 191 120 208
rect 328 207 345 224
rect 205 170 222 187
rect -35 121 -18 138
rect 430 248 447 265
rect 509 207 526 224
rect 274 143 291 160
rect -191 87 -169 109
<< metal1 >>
rect 104 306 345 320
rect 104 264 120 306
rect -239 250 120 264
rect -239 232 -222 250
rect -247 224 -214 232
rect -247 207 -239 224
rect -222 207 -214 224
rect -247 199 -214 207
rect -93 224 -60 232
rect -93 207 -85 224
rect -68 207 -60 224
rect -93 199 -60 207
rect 19 215 52 223
rect 103 216 120 250
rect 328 232 345 306
rect 371 306 404 315
rect 371 289 378 306
rect 396 289 526 306
rect 371 281 404 289
rect 422 265 455 273
rect 422 248 430 265
rect 447 248 455 265
rect 422 240 455 248
rect 320 224 353 232
rect -86 176 -69 199
rect 19 198 27 215
rect 44 198 52 215
rect 19 190 52 198
rect 95 208 128 216
rect 95 191 103 208
rect 120 191 128 208
rect 320 207 328 224
rect 345 207 353 224
rect 320 199 353 207
rect 29 176 46 190
rect 95 183 128 191
rect 197 187 230 195
rect -239 162 46 176
rect 197 170 205 187
rect 222 170 230 187
rect 197 162 230 170
rect -239 54 -225 162
rect -42 142 -9 143
rect 205 142 222 162
rect -42 138 222 142
rect -42 121 -35 138
rect -18 127 222 138
rect 266 160 299 168
rect 266 143 274 160
rect 291 143 299 160
rect 266 135 299 143
rect -18 121 -9 127
rect -42 115 -9 121
rect -196 109 -163 115
rect -196 87 -191 109
rect -169 88 -163 109
rect 274 88 291 135
rect -169 87 291 88
rect -196 72 291 87
rect 430 54 450 240
rect 509 232 526 289
rect 501 224 534 232
rect 501 207 509 224
rect 526 207 534 224
rect 501 199 534 207
rect -239 40 450 54
use inv  inv_0
timestamp 1679616770
transform 1 0 502 0 1 62
box -42 -62 121 426
use inv  inv_1
timestamp 1679616770
transform 1 0 -92 0 1 62
box -42 -62 121 426
use inv  inv_2
timestamp 1679616770
transform 1 0 -246 0 1 62
box -42 -62 121 426
use nand2  nand2_0
timestamp 1676660346
transform 1 0 321 0 1 62
box -42 -62 175 426
use xor2  xor2_0
timestamp 1677800174
transform 1 0 42 0 1 62
box -42 -62 283 426
<< labels >>
flabel locali s -93 199 -60 232 0 FreeSerif 80 0 0 0 B
port 2 nsew
flabel locali s -247 199 -214 232 0 FreeSerif 80 0 0 0 A
port 1 nsew
flabel locali s 200 216 233 281 0 FreeSerif 80 0 0 0 S
port 0 nsew
flabel locali s 552 115 585 315 0 FreeSerif 80 0 0 0 C_out
port 6 nsew
flabel locali -286 432 621 480 0 FreeSerif 80 0 0 0 VDD!
flabel locali s -286 0 621 48 0 FreeSerif 80 0 0 0 GND!
<< end >>
