magic
tech sky130A
magscale 1 2
timestamp 1681866284
<< locali >>
rect -264 864 3238 960
rect -84 331 -18 630
rect 82 528 148 594
rect 1654 528 1720 594
rect 286 483 484 494
rect 286 449 373 483
rect 407 449 484 483
rect 286 428 484 449
rect 1858 477 2056 494
rect 1858 443 1941 477
rect 1975 443 2056 477
rect 1858 428 2056 443
rect -84 265 -62 331
rect -84 230 -18 265
rect 1164 261 1230 394
rect 1500 230 1566 394
rect 2736 230 2802 394
rect 3072 230 3138 394
rect 1183 226 1211 227
rect -264 0 3238 96
<< viali >>
rect -186 398 -120 464
rect 373 449 407 483
rect 1941 443 1975 477
rect -62 265 -18 331
rect 1164 227 1230 261
<< metal1 >>
rect 361 488 419 489
rect 27 483 419 488
rect -192 464 -114 476
rect -192 398 -186 464
rect -120 454 -114 464
rect 27 454 373 483
rect -120 449 373 454
rect 407 449 419 483
rect -120 443 419 449
rect -120 409 72 443
rect -120 398 -114 409
rect -192 386 -114 398
rect -68 331 -12 343
rect -68 265 -62 331
rect -18 318 -12 331
rect -18 278 180 318
rect -18 265 -12 278
rect -68 253 -12 265
rect 140 163 180 278
rect 1152 261 1242 267
rect 1152 227 1164 261
rect 1230 258 1242 261
rect 1678 258 1706 578
rect 1929 478 1987 483
rect 1230 230 1706 258
rect 1763 477 1987 478
rect 1763 443 1941 477
rect 1975 443 1987 477
rect 1763 441 1987 443
rect 1230 227 1242 230
rect 1152 221 1242 227
rect 1763 163 1800 441
rect 1929 437 1987 441
rect 140 126 1800 163
rect 140 124 180 126
use Dlatch  Dlatch_0
timestamp 1679435600
transform 1 0 84 0 1 124
box -84 -124 1586 852
use Dlatch  Dlatch_1
timestamp 1679435600
transform 1 0 1656 0 1 124
box -84 -124 1586 852
use inv  inv_0
timestamp 1679616770
transform 1 0 -184 0 1 124
box -84 -124 242 852
<< labels >>
flabel locali s -186 398 -120 464 0 FreeSerif 400 0 0 0 CLK
port 5 nsew
flabel locali s 82 528 148 594 0 FreeSerif 400 0 0 0 D
port 0 nsew
flabel locali s 2736 230 2802 394 0 FreeSerif 400 0 0 0 Q
port 1 nsew
flabel locali s 3072 230 3138 394 0 FreeSerif 400 0 0 0 NOT_Q
port 2 nsew
<< end >>
